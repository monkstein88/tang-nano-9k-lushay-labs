// In this article we will be taking a look at generating pseudo-random numbers using an LFSR (Linear Feedback Shift Register) and look at how one can be used as part of a larger application.
//
// The LFSR
// An LFSR is a shift register like we have seen in previous articles, except that the bits besides shifting are also affected by the other bits in the register - this effect is what is referred 
// to as the feedback.
//
// There are multiple variations of LFSR but in this article we will be focusing on the most basic type the Fibonacci LFSR. In this type of LFSR the feedback only affects the first bit. So all 
// bits get shifted up and the least significant bit is generated using the feedback of the current registers bits.
// 
// A basic example of a 5-bit LFSR:
//
//                                /-----|| 
//                               /      ||<----------------------+
//               +--------------{  XOR  ||                       |
//               |               \      ||<--+                   |
//               |                \-----||   |                   |
//               |                           |                   |
//               |                           |                   |
//               |                 +-----+---*--+------+-----+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |  B3 |  B4  |-------| >
//                 LSFR INPUT BIT  |     |      |      |     |      |       |/
//                                 +-----+------+------+-----+------+
//                                   LSb                        MSb
//                                     
// So in the example above on each clock cycle B4 is the output bit b0-b3 get shifted up and a new bit is generated by XOR-ing bit 4 and bit 1 this new bit gets inserted into b0.
//
// The bits we choose for our feedback are called "taps", and not every arrangement of taps are good options. Since our new bit is generated by XOR-ing bits, if all bits were zero the system 
// would be stuck in the zero state. XOR can be thought of as returning 1 if the number of 1s being XOR-ed is odd. Since all zeroes has zero 1s and shifting will just keep inputting a new zero
// we never get out of this state.
//
// Another thing to consider, the entire equation is only based on the current state of the register there is no other state being used in the calculation, so as soon as the register rolls 
// back to a number it already was on that will create a cycle. For example if we have an LFSR generating numbers from 1-16 but has an initial cycle of: 1, 4, 7, 14, 3, 5, 7, 14, 3, 5, 7
//
// You can see that as soon as we had two ways of getting to 7 (both 4 generated a 7 as the next number and also a 5) we get stuck in a loop between the two numbers. All further cycles will just
// go between 7, 14, 3, 5 in an endless cycle.
//
// The problem with these short cycles is that the LFSR can no longer generate any number in the range. If I have a 6-sided dice that can only be a 2 or a 4 it wouldn't really be considered a 
// fair dice in the realm of numbers 1-6 as the probabilities for each number are not the same.
//
// So when choosing taps we want to choose something that:
// 1. Never generates all zeroes
// 2. Generates a sequence that goes through all possible numbers
//
// Luckily for us, we do not have to manually calculate optimal taps instead there are pre-calculated tables for max length taps. For example this site here has a precompiled list of max-length 
// taps for LFSRs with 4-64 bits.
//
// For example opening the file for 5-bit LFSRs like in the example above has the following options:
// 0x12
// 0x14
// 0x17
// 0x1B
// 0x1D
// 0x1E
//
// Each of these is an optional tap set. The example above used the 12 option, these numbers are in hex, but converting 12 hex to binary provides:
// 0b10010
//
// Least significant bit to least significant bit, this means take bits index 1 and index 4 for the feedback and leave out index 0,2 and 3 like in this image:
//
//                                /-----|| 
//                               /      ||<----------------------+
//               +--------------{  XOR  ||                       |
//               |               \      ||<--+                   |
//               |                \-----||   |                   |
//               |                           |                   |
//               |                           |                   |
//               |                 +-----+---*--+------+-----+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |  B3 |  B4  |-------| >
//                 LSFR INPUT BIT  |     |      |      |     |      |       |/
//                                 +-----+------+------+-----+------+
//                                   LSb                        MSb
//
// But any of these options would produce a max-length sequence. Now that we have something that can generate a complete sequence of all numbers let us talk a little about the "random" part.
//
//
// Pseudo Random
//
// The LFSR produces a sequence which includes all the possible options, but that doesn't necessarily make it "random". For example if we are talking about a 3-bit LFSR, we can get all the numbers
// 1-7, but a 3-bit counter also produces all the numbers from 1-7 but it would hardly be random.
//
// Taking a look at a counter's sequence:  
// 1,2,3,4,5,6,7
//
// All numbers in this sequence have the same number of occurrences, but each number is just the previous number plus 1 making it to obvious of a relationship for us to call it unpredictable 
// or random.
//
// Now like with a deck of cards, the way can randomize the output is by shuffling. So let's shuffle this group of numbers into the following for example:
// 7, 6, 4, 1, 2, 5, 3
//
// One can now say that the sequence is random, because the order in which the numbers come out are no longer related to previous elements. The sequence is still not perfect as there are no duplicates,
// for example with rolling a dice I can roll a 4 and then roll another 4 before going through all the other options. But we can at least say it is as random as a deck of cards being randomly shuffled.
// 
// The problem with this solution is it requires something else to randomly shuffle the elements for it to really be random and it is hardware intensive to implement. To create such a system we would 
// need to store each number of the sequence kind of like a 1-time pad so for example with a 32-bit LFSR we would need to store 2^32 -1 numbers over 4-billion 32-bit numbers or about 16GB of storage 
// for 1 sequence, and we would even want sequences much longer then this.
//
// So an LFSR is somewhere in-between a real shuffled sequence to a sequence with an obvious relation like a counter. The LFSR - when the taps are chosen correctly - produces all the numbers (except 0)
// in a sequence shuffled based on a non-obvious relation.
//
//
//                                /-----||      
//                               /      ||<---------+
//               +--------------{  XOR  ||          |
//               |               \      ||<--+      |
//               |                \-----||   |      |
//               |                           |      |
//               |                           |      |
//               |                 +-----+---*--+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |-------| >
//                 LSFR INPUT BIT  |     |      |      |       |/
//                                 +-----+------+------+
//                                   LSb           MSb
//
// Starting with the seed value (initial value) of 1, let's the sequence given by this shift register will be:
// binary  | decimal
//  001    | 1
//  011    | 3
//  111    | 7
//  110    | 6
//  101    | 5
//  010    | 2
//  100    | 4
//  001    | 1
//
// Looking at this sequence you can see that we go through all the numbers before reaching back to 1 and that the sequence is shuffled. The reason we call this "pseudo-random" and not random is because 
// there is a correlation between them, it can be said that the function for the first bit is:
// b0 = b1 xor b2
// and that for the other bits the equation is simply:
// b_i = b_(i-1)
//
// As each bit is simply shifted up. Since there is a correlation between the previous state and the next state with enough of the sequences outputs one could solve some math equations and work out which 
// taps were chosen being able to predict future numbers in the sequence.
//
// So it's not unpredictable, but the order has no meaningful meaning so we can say it is shuffled. With that said there are some things we can do to make it even better.
//
// The first thing is to make the LFSR larger then the number we are using. For example if we need a 4-bit number and we use instead a 5-bit LFSR taking 4 bits at a time, we essentially doubled the number
// of times each number comes up allowing our sequence to have streaks of the same number like we mentioned that dice rolls have. We also get the ability to get 0 as a number, all the bits of an LFSR 
// cannot equal zero but if you are reading only some of the bits then they can all equal zero.
//
// In reality you usually want the LFSR to be much bigger (not just by one bit) and use a relatively small number of bits. Another way to make it better is to not reuse the same bits and to skip bits 
// in-between numbers.
//
// Each shift of the register you only get 1 new "random" bit. All the other bits are just shifted over which is like doubling. So in the case of the 3-bit LFSR if you wait 3-bits before taking another
// number then all of the new numbers 3-bits are completely unrelated to the bits of the previous number making it more random.
//
// Finally if you let the LFSR run in the background essentially skipping generated bits and then let random actions like when a user pressed a button decide when to read the next number you are 
// essentially adding in random like when shuffling bringing it closer to real random.
//
// I think that is enough theory though let's get into building this.
//


module top
#(
  /* Tang Nano 9K Board - featuring GOWIN FPGA: GW1NR-LV9 QFN88P (rev.C) */
  parameter EXT_CLK_FREQ = 27000000, // external clock source, frequency in [Hz], 
  parameter EXT_CLK_PERIOD = 37.037, // external clock source, period in [ns], 
  parameter STARTUP_WAIT_MS = 10 // make startup delay of 10 [ms]
)
(
  input wire EXT_CLK,  // This is the external clock source on the board - expected 27 [MHz] oscillator. 
  input wire BTN_S1, // This pin is tied to a button 'S1' on the board, and will be used as a 'reset' source (active-low) 
  input wire BTN_S2, // This pin is tied to a button 'S2' on the board, and will be used as a general user input source (active-low) 
  output reg [5:0] LED_O=6'b1, // 6 Orange LEDs on the board, active-low , default to all high (leds are OFF)
  // LCD 0.96" SPI interface - SSD1306 controller
  output wire LCD_RST, // reset: active-low   
  output wire LCD_SPI_CS, // chip-select: active-low Note: multiple bytes can be sent without needing to change the chip select each time.
  output wire LCD_SPI_SCLK, // spi clock signal: idle-low 
  output wire LCD_SPI_DIN, // data input. Note: data is latched on the rising edge of the clock and is updated on the falling edge. MSb is sent first.
  output wire LCD_DC,  // data/command select: active-low - data, active-high - command

  input  wire UART_RX, // UART|RX pin - 8N1 config
  output wire UART_TX,  // UART|TX pin - 8N1 config
  
  output wire FLASH_SPI_CS,  // chip select for flash memory
  output wire FLASH_SPI_MOSI, // master out slave in for flash memory
  input  wire FLASH_SPI_MISO, // master in slave out for flash memory
  output wire FLASH_SPI_CLK  //  clock signal for flash memory
);
localparam STARTUP_WAIT_CYCL = ((EXT_CLK_FREQ/1000)*STARTUP_WAIT_MS);

wire  [9:0] pixelAddress;
wire  [7:0] textPixelData;

// Let's now take a look if we don't reuse bits and only take 3-bit numbers.
wire randomBit; // creating a wire for the randomBit
lfsrTest testLFSR( // creating an instance of our test LFSR connecting it to our wire.
  clk,
  randomBit
);
reg [2:0] tempBuffer = 0; // create a buffer to hold the bits as they are shifted off the LFSR
reg [1:0] counter = 0; // create another register to count every time we got 3 new bits 
reg [2:0] value; // and a final register to store the value once ready.

always_ff @(posedge clk) begin  // Inside the clock loop ...
  if(counter == 3) begin  // ... we check for when the counter reaches 3 ... 
    value <= tempBuffer; // ...  in which case we transfer the temp value into the value register.
  end
  counter <= counter + 1; // Other then that we always increment the counter ... 
  tempBuffer <= {tempBuffer[1:0], randomBit}; // ...  and shift the new randomBit into our temp buffer shifting everything up.
end
// Looking at the output of this - The first two numbers are not defined ('z') as we didn't initialize our registers with a value but it's ok since not all the bits are random there.
// Looking at the sequence now we get: 2,3,3,1,7,3,4,0,5,7,6,3,6,6,1,0,2,6,4,7,4,5,2,1,5,5,0,7,1,2,4
//
// Our sequence length is still 31 but now since we are reading smaller bit-sized numbers we have multiple duplicates of each number 4 to be exact since we left off two bits and 2^2 = 4.
// Except for 0 which there is only 3 since one of the options is when the LFSR equals all zeros which is not a valid case.
//
// Another benefit here is you can see there are some streaks and also if you get a number for example a 2 you don't know the next number as it could be a 3,6,1 or 4 because of the multiple occurrences.
//
// Adding the fact that you let it run at 27MHZ that means it goes through the whole cycle about 900,000 times a second or about 1 micro-second. If you only take a number based on for example user-input
// like a button press, a person can't reliably time their button presses to 1/31-th of a microsecond to get a specific number in the sequence making it pretty much random for most use-cases.
//
// Before we start playing with LFSRs let's see how we can generalize our module so we don't need to create a new one for each different LFSR we add.
endmodule

// The Implementation
// Implementation wise it couldn't be any easier we just need a register with the number of bits we want in the LFSR and we need to connect some of the bits to the input of the first bit based on 
// the taps we chose.
// 
// Taking our 5 bit LFSR from before we can create a simple verilog file like the following:
module lfsrTest(
  input   wire  clk, 
  output   reg  randomBit = 0
);

  reg  [4:0] sr = 5'b00001;
  
  always_ff @(posedge clk) begin 
    sr <= {sr[3:0], sr[4] ^ sr[1]};
    randomBit <= sr[4];
  end
// We seed the shift register with an initial value of 1 and on each clock pulse we shift the bits up and calculate the new input bit for b0 by XOR-ing bit 4 and bit 1 together. We then set the output 
// register which holds the random bit to the value of b4 in our shift register (the bit we shifted off).
// 
// Running this would produce the following sequence:
// 1,2,5,10,21,11,23,14,29,27,22,12,24,17,3,7,15,31,30,28,25,19,6,13,26,20,9,18,4,8,16
//
// With five bits we have 2^5 options -1 removing the zero case we get a period of 31 numbers. And as you can see the order seems pretty random. Already looks pretty good but again there is some
// correlations where you can see the number just doubling because of the shift for example at the beginning or end of the sequence.
endmodule