//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.03 (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Aug 17 00:03:07 2025

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din);

output [3:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [15:0] ad;
input [3:0] din;

wire lut_f_0;
wire [30:0] sp_inst_0_dout_w;
wire [0:0] sp_inst_0_dout;
wire [30:0] sp_inst_1_dout_w;
wire [0:0] sp_inst_1_dout;
wire [30:0] sp_inst_2_dout_w;
wire [1:1] sp_inst_2_dout;
wire [30:0] sp_inst_3_dout_w;
wire [1:1] sp_inst_3_dout;
wire [30:0] sp_inst_4_dout_w;
wire [2:2] sp_inst_4_dout;
wire [30:0] sp_inst_5_dout_w;
wire [2:2] sp_inst_5_dout;
wire [30:0] sp_inst_6_dout_w;
wire [3:3] sp_inst_6_dout;
wire [30:0] sp_inst_7_dout_w;
wire [3:3] sp_inst_7_dout;
wire [30:0] sp_inst_8_dout_w;
wire [0:0] sp_inst_8_dout;
wire [30:0] sp_inst_9_dout_w;
wire [1:1] sp_inst_9_dout;
wire [30:0] sp_inst_10_dout_w;
wire [2:2] sp_inst_10_dout;
wire [30:0] sp_inst_11_dout_w;
wire [3:3] sp_inst_11_dout;
wire [29:0] sp_inst_12_dout_w;
wire [1:0] sp_inst_12_dout;
wire [29:0] sp_inst_13_dout_w;
wire [3:2] sp_inst_13_dout;
wire [27:0] sp_inst_14_dout_w;
wire [3:0] sp_inst_14_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_44;
wire mux_o_45;
wire mux_o_46;
wire ce_w;
wire gw_gnd;

assign ce_w = ~wre & ce;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[12]),
  .I1(ad[13]),
  .I2(ad[14]),
  .I3(ad[15])
);
defparam lut_inst_0.INIT = 16'h4000;
SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[30:0],sp_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 1;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hFFEFFDEFFFFFFFFFFFFFFFFFDC7FFEFDFFF4340000005FDB823FFEFFFFFF91FF;
defparam sp_inst_0.INIT_RAM_01 = 256'hFFDDF7FFEFFFFFFFFFFFFFFFF5EFFFFDF5DA025020407BF6DF3FFFFFFFFD0AFF;
defparam sp_inst_0.INIT_RAM_02 = 256'hFFD5F57FFFFFEFFFFFFFFFFFF77FEFBFF6D34901C3011E5E08DFFFFFFFFC10FF;
defparam sp_inst_0.INIT_RAM_03 = 256'hFCBDFFFFFFFFFFFFFFFFFFFFFFFDFFB5FFEEFE25801565907A1FFFFFFCBC14FF;
defparam sp_inst_0.INIT_RAM_04 = 256'hF05C5FFFFFDFFFFFFFFFFFFFFFFFAFFF6FDFFF7DC0C5FBC59C5FFFFFFBDE403F;
defparam sp_inst_0.INIT_RAM_05 = 256'hC0FFFFBFFFFFFFFFFFFFFFFFFFFFFFFF3FFBED9BE02EFB152EC7FFFFFEB0020F;
defparam sp_inst_0.INIT_RAM_06 = 256'h00CFF76FFFFFFFFFFFFFFFFFFFDFFFF3FDF3DFFB733DE91CD8BFFFFDFFA00003;
defparam sp_inst_0.INIT_RAM_07 = 256'h00FFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBBFBABD11AC76FFFFFFC200000;
defparam sp_inst_0.INIT_RAM_08 = 256'h00D9EDFFDFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFBFFF42A7AFFFFFFD800000;
defparam sp_inst_0.INIT_RAM_09 = 256'h00FFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBFFE180097BF7FFB4000000;
defparam sp_inst_0.INIT_RAM_0A = 256'h00BFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF7FFFF25E299EBFFFE38000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFBF1CE9E7FE7F64000000;
defparam sp_inst_0.INIT_RAM_0C = 256'h00FDBFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFDF5F4481BFDF000000000;
defparam sp_inst_0.INIT_RAM_0D = 256'h00FFFBFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFF7FFFFFCA9051006F76301000000;
defparam sp_inst_0.INIT_RAM_0E = 256'h00FDEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFF996B259F1EE1000000400;
defparam sp_inst_0.INIT_RAM_0F = 256'h00FFEFFFFFFFF7FFFFFFEFFFFFFFFFFFFFFFFFFBFFF58A01D17BF20000000000;
defparam sp_inst_0.INIT_RAM_10 = 256'h00F5FFFFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFF347830701FDA000000000;
defparam sp_inst_0.INIT_RAM_11 = 256'h00BFFFFFFFFFFEFEFFFFFFFFFFFFFFFFFFFFFFB7FFF7A67714EFFE0820000000;
defparam sp_inst_0.INIT_RAM_12 = 256'h00EFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFCA2A2AEA37FDA000000000;
defparam sp_inst_0.INIT_RAM_13 = 256'h01FFFFF7DFFFFDFFFF7FFFFFFFFFFFFFFFFFFFFFFFE04DC0BFBBF70000000000;
defparam sp_inst_0.INIT_RAM_14 = 256'h07FFFFFDFFFFFFFEFFFFFFFFFFFFDFFFFFFFFFFFFFDCCB5638A3F5A000000080;
defparam sp_inst_0.INIT_RAM_15 = 256'h1FFFFFFFFFFFFFFFDF9FFFFFFFFFFFFFFFFFFFFFFF99C719ECF6FE01000000E0;
defparam sp_inst_0.INIT_RAM_16 = 256'h7FFFDBEFFFFFFFFF7FFFFBFFFFEFFFFFFFFFFFFFFFE6AEDA675A98B0000000F8;
defparam sp_inst_0.INIT_RAM_17 = 256'hFFFFB7FFFFFCFFBFFFEFDFFFFFFFFFFFFFFFFFFFEE07EB9F01D7EA10000000FE;
defparam sp_inst_0.INIT_RAM_18 = 256'hFFFFD7DF7FBFFFBFFFFFFFFFFFFFFFFDFFFFFFFFFF61C7ECA9BECC00000000FF;
defparam sp_inst_0.INIT_RAM_19 = 256'hFFFFEFFFBDFFDFDFF3BFDFFFFFFFFFFFFFFFFFFFFE431A96FC753000000000FF;
defparam sp_inst_0.INIT_RAM_1A = 256'hFFFFF7DFFF3FFFFFFE6FFFFFFFFFFFFFFFFFFFFFFAEAEB51E023A000000000FF;
defparam sp_inst_0.INIT_RAM_1B = 256'hFFFAFBFFF95BFFEFBFFFEFFFFFFFFFFFFFFFFFFFFEE73D823587E000000000FF;
defparam sp_inst_0.INIT_RAM_1C = 256'hFF7FF6DF7FBFEAFFFFFFFFDFFFFFFFFFFFFFFFFFE6B2F2069216C000000000FF;
defparam sp_inst_0.INIT_RAM_1D = 256'hFFF7CFFFFDD7FEFFFFFFDFFFFFFFFFFFFFFFFFFFEF9C8720045F0000000000FF;
defparam sp_inst_0.INIT_RAM_1E = 256'hFFF67D7E77DFEFFFFFFFFFFFFFFFFFFFFFFFFFFFCC0F9EEBE2B3C000000000FF;
defparam sp_inst_0.INIT_RAM_1F = 256'hFFFF3FFFF76FBFFFFDFEFFFFFFFFFFFFFFFFF3FFDF0ACBD1CD8F0000000001FF;
defparam sp_inst_0.INIT_RAM_20 = 256'hFFDDDAFFFF7FFD7FEFFFF7FFFFFFFFFFFFDFFFFFB5309DCE8B6C0000000000FF;
defparam sp_inst_0.INIT_RAM_21 = 256'hFF6B0FFE7BFF7FDFFFFFFFFFFFFFFFFFDFFDD6FB73673205E8D40000000002FF;
defparam sp_inst_0.INIT_RAM_22 = 256'hFF7E1CBA7EB3FBFFFFFEFFFFFFFFFFFFFFFDDBFED05B691E7BE7D800000000FF;
defparam sp_inst_0.INIT_RAM_23 = 256'hFFA766C9EEF8ABFFFFFFFFFFFFFFFFFFFFFBBBDED353B3807E4E3000000000FF;
defparam sp_inst_0.INIT_RAM_24 = 256'hFF947DB77EF7FFFFFF9FFFFFFFFFFFFFBFFFB389B35AD7E088378000000040FF;
defparam sp_inst_0.INIT_RAM_25 = 256'hFCC0759AC7DFFFFFFFFF7FFFFFFFDEFF7FFFEAE3E6ACC890B3C59000000043FF;
defparam sp_inst_0.INIT_RAM_26 = 256'hF06B1ED337EFFFFFFFFFFFFFFFFFFFFFFFFD10A4291BACFE439C000000001A3F;
defparam sp_inst_0.INIT_RAM_27 = 256'hC06D38643BEEFFFFFFFFFFFFFFFFFFFFFDF77B2BFDFE2C60A26300000000000F;
defparam sp_inst_0.INIT_RAM_28 = 256'h00208A2C4F1FFFFDFFFDFFFFFFFFFCFFFFBFE3EDF4D31C67C066000000008C03;
defparam sp_inst_0.INIT_RAM_29 = 256'h00888928DDFFEFFFB7FEFFFBFFFFFFFFF6CAE28DB22FFC70C3CE000000000100;
defparam sp_inst_0.INIT_RAM_2A = 256'h00BB06AA6EE5FFFFFFFFFFFFFFFFFDFFFFE1F11BE41DDF7834C4000000004100;
defparam sp_inst_0.INIT_RAM_2B = 256'h001000553012FFFDFFFF7FFFFFFFFFFFEDFA280BEE7791DF8BC8600000408000;
defparam sp_inst_0.INIT_RAM_2C = 256'h0008110B71BF7DDF7DFFFFFFFFFFFFFFDF93A023EF7AF65B2046F00000200100;
defparam sp_inst_0.INIT_RAM_2D = 256'h00006007EFCCFF3EBBFFFFFFFFFFFFFFFFB7C051C11A4AA0A213A80008047400;
defparam sp_inst_0.INIT_RAM_2E = 256'h003A7C9CF4D57FFEFFFFFFFFFFFFFFFFFBDFE04DCAB888E30110FE0000020000;
defparam sp_inst_0.INIT_RAM_2F = 256'h006D5A9CFAF3FFFFFFFFFFDFFFFFFBFFDFDFC4D3C7F908009410A80000880100;
defparam sp_inst_0.INIT_RAM_30 = 256'h00413BB1BC4BBFF7FFFFFFFFFDFFFDFDFFDFC607EDCE04491FFE380802800000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0012CE80ABFEFFFFFFFFDFBFFFFFFF7DFBDF8EA5EFCB42E4FF44000000A70400;
defparam sp_inst_0.INIT_RAM_32 = 256'h005B65ED2596FFDFFFFFFFFFBFFFFFBD77DC0697C74A6FDC5FBC800000290100;
defparam sp_inst_0.INIT_RAM_33 = 256'h00066E18D07EF2F7FFFFBEF7DFFFFFFEFBCA05DFA659A7FE0F3D7A0000D12000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0067F0706D49DFFDFF7FFBFFFFFFFFFFEC205837C749F7DD6E75800000802900;
defparam sp_inst_0.INIT_RAM_35 = 256'h01663221CDE137FFFFFFFDFD76FFFFFC0441059FEC43F1C87FDA500000783400;
defparam sp_inst_0.INIT_RAM_36 = 256'h07EBA3303D5C3BFBFFFFFFFFFFFFFFEC000206EFF90CA0F88FC3B00000011680;
defparam sp_inst_0.INIT_RAM_37 = 256'h1FBB9F999C40BFFFFFFFFFFFEBFFFC6002C41DF9F188BF89F80010020C1204E0;
defparam sp_inst_0.INIT_RAM_38 = 256'h7F1FF0303F006FDF7FFFDF9FE7FFC4281A494A3F4303FE703C0E0080400080F8;
defparam sp_inst_0.INIT_RAM_39 = 256'hFF9FD3FF33CE2E7FFFF7FFFFFFFD2428201892FF9B638967F80A0001868285FE;
defparam sp_inst_0.INIT_RAM_3A = 256'hFFFF1FF7AAA7ECFFFFFFFFBFEFB0003004FFC35F1681F113F916000001330EFF;
defparam sp_inst_0.INIT_RAM_3B = 256'hFF6D3E679FE9AEEDFFFFFFFFCF8000890DFFF3E54B340051F8D8000122007CFF;
defparam sp_inst_0.INIT_RAM_3C = 256'hFFF8BE7E0930FBFF7FFFFFFFFC000CE41BFFE7F69307B7B8F1EA0000000388FF;
defparam sp_inst_0.INIT_RAM_3D = 256'hFFE957E495FF05F7FBEFFDFAF62402586417F6B6E9CC7350706F00000006F9FF;
defparam sp_inst_0.INIT_RAM_3E = 256'hFFB18078E8F2B9AFFFFEF8A02033C8B4DB02E7D84708C337B00D0000010342FF;
defparam sp_inst_0.INIT_RAM_3F = 256'hFFBE10DB3A03162AF7FFDA0080022580FCDCFF8F50E8676301E280000865E3FF;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[30:0],sp_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 1;
defparam sp_inst_1.BLK_SEL = 3'b001;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'hFF742B15D802E751BFFFD40604814FC9FFCDD7FE716E0B2487F3A000000883FF;
defparam sp_inst_1.INIT_RAM_01 = 256'hFFF83202901382062B9BE06E8E490FE5FF331CDC39A4CC31FF7BB000001051FF;
defparam sp_inst_1.INIT_RAM_02 = 256'hFF181D8374166151038BF0FF1AD80F80F06C27DC3143BF50FBF91000010806FF;
defparam sp_inst_1.INIT_RAM_03 = 256'hFF3811F7CEFA782B4043F86FB0F90FFBFC9C69ECAA6E73A1F3FA3000054211FF;
defparam sp_inst_1.INIT_RAM_04 = 256'hFF31695832F503FDF030056BFBFF0703244E6ECA64F827C72FF53010024E62FF;
defparam sp_inst_1.INIT_RAM_05 = 256'hFF24BD8A1383A03D44AA97032BFF27F7FC4A87EDD53EECE356E9800016095FFF;
defparam sp_inst_1.INIT_RAM_06 = 256'hFF05DD23775E11C35980E73F8BFE0782FC3EC14E5FF01133E1E8200001A985FF;
defparam sp_inst_1.INIT_RAM_07 = 256'hFCB86D163B647233A9929B8BC1FA07AF967A2F685F32B762C7A600000C7506FF;
defparam sp_inst_1.INIT_RAM_08 = 256'hF0D75DAC15151A1F1149EFEDC8E3079E4C414F269CBDDFD0FB8CE0000199183F;
defparam sp_inst_1.INIT_RAM_09 = 256'hC0CB1DACB60A70CAF9D73FEF60EB83C60B486A5AF3A43B7193B2D0010642100F;
defparam sp_inst_1.INIT_RAM_0A = 256'h00AF0B91AE117E5ED956FB7CC2A7DFC00DE7B952D76BED68819B400005CE3403;
defparam sp_inst_1.INIT_RAM_0B = 256'h0068787C1D635F83FD0FFDD903AFBB84C7587E0971C193BC686D140010B30400;
defparam sp_inst_1.INIT_RAM_0C = 256'h001A9F53043DE3D0FF157FD96B33C3B1E612EB5644B7FAEFF62EF00001842A00;
defparam sp_inst_1.INIT_RAM_0D = 256'h007BBF4F5A23FC947E357260DFE9E1F1094FFDDDBE7EB45921E63000108A1200;
defparam sp_inst_1.INIT_RAM_0E = 256'h00BB8772C6EB5FF3D9F8E001EB05ADEAD62D8F9E02D694769E61800072559D00;
defparam sp_inst_1.INIT_RAM_0F = 256'h0041E177093B0BD06DFFE1B191E7EFAA2B88E5D61C0D86249E68300001208B00;
defparam sp_inst_1.INIT_RAM_10 = 256'h006C8BFB9AE300FCBF7E96B1A3A5E7CDCAC097B76E57508005FE500004B14C00;
defparam sp_inst_1.INIT_RAM_11 = 256'h00EAA76F35E188885EFFD7C1FB595FC381C8CBBDAF7BF28B67FDB000020C9700;
defparam sp_inst_1.INIT_RAM_12 = 256'h000580A40ABFDEFE3F7D45A4FBC79F55E7F435E9797AB8BF2FFFA00081680000;
defparam sp_inst_1.INIT_RAM_13 = 256'h002F6CD01F7D6498CD7F5BC2F3060E96AB90202691F960D32DAA04002B840000;
defparam sp_inst_1.INIT_RAM_14 = 256'h00E5C92C26EE9DBC53BE918FAFD0A397FBF466EEE18FB43D5DB406000E200000;
defparam sp_inst_1.INIT_RAM_15 = 256'h002223503EDFDDE2A6CFEF0783F2E9FE5A7B7EBB39FBCD1799C0010052B50000;
defparam sp_inst_1.INIT_RAM_16 = 256'h00539B87B9075FD85BFBAE8FA559EBB3C1ECF13F97BEDBAA69294E02CBF00900;
defparam sp_inst_1.INIT_RAM_17 = 256'h01106FE539A35C0F6348ED8EE0B2701E7D61F3CD97EBCFE66AE0050000B10900;
defparam sp_inst_1.INIT_RAM_18 = 256'h07002BB6F598EE0D46DBFC9BD8B26CAD7E97AA1744DB668FC8C97F4002500580;
defparam sp_inst_1.INIT_RAM_19 = 256'h1F893D3D76B930A972CBF91E93DD2C7995D2B528EE15FBB473B23EA2009000E0;
defparam sp_inst_1.INIT_RAM_1A = 256'h7F8724F3172E70E6CF8FFAF9C641CF0F046394A10C457A3195F0F4B005A004F8;
defparam sp_inst_1.INIT_RAM_1B = 256'hFF0698C0B87117C049BF1C988F17FEBD061DEF64A84522BEA3F89DA000DC06FE;
defparam sp_inst_1.INIT_RAM_1C = 256'hFF0428D4A5CEAC17A37FEF24BC477C19868F1941D644DAD706C0FA00203206FF;
defparam sp_inst_1.INIT_RAM_1D = 256'hFF043D27066191203354A44B7EEDF7A0814454C5A80677C4F470F2B9000000FF;
defparam sp_inst_1.INIT_RAM_1E = 256'hFF08E04912C7AEF9A0367CBAD662F7D84A2F966B6C9FB95A95CCFB6A008000FF;
defparam sp_inst_1.INIT_RAM_1F = 256'hFF16002A898267A48BFC92A76DD1FFAB8C380CF1600F1D5FA715A342000000FF;
defparam sp_inst_1.INIT_RAM_20 = 256'hFF0E5BCC3729B54DFFE80CEA4A7EF711D16607A9803721FA64068AD2800040FF;
defparam sp_inst_1.INIT_RAM_21 = 256'hFF01CDE44B9B115D2DD5043A69B9F96A1FC347E185635EF80A5791FE002E19FF;
defparam sp_inst_1.INIT_RAM_22 = 256'hFF008227A822C6F8CF9FFEFB12C2FD6F0C5A83F6DBE9A7416B2BC9F8819C6FFF;
defparam sp_inst_1.INIT_RAM_23 = 256'hFF000259558240D517EB56C3725CA8C20D5BA0ED4D41FE969C93A9C0C773A3FF;
defparam sp_inst_1.INIT_RAM_24 = 256'hFF001017982F811DD0B5D0FEEC5D12330009A0FC0E38B327A0F63A3C7F7F43FF;
defparam sp_inst_1.INIT_RAM_25 = 256'hFF0006BF3C171A33EDFC42F5B435DE3FB27530CE55E32503CF9F277C7F081BFF;
defparam sp_inst_1.INIT_RAM_26 = 256'hFF000A93B86FFABC4201A79EAA0EAE711C64B01CAA4ADA94B816B8361FE83FFF;
defparam sp_inst_1.INIT_RAM_27 = 256'hFF010EB7C00EFFB30D28B656781B7A7D1991588D210E4E8E6AA1D54C13F93FFF;
defparam sp_inst_1.INIT_RAM_28 = 256'hFF020D1D6FFD9326FA1EFAFDB60AB51300CADDEBEFE62562CEBEA6109BF05FFF;
defparam sp_inst_1.INIT_RAM_29 = 256'hFC0008F0170A41A466D0B172E0027F890C2D96768BDCC40BFBB64FC30F38C8FF;
defparam sp_inst_1.INIT_RAM_2A = 256'hF0000E584725D38024B1617A080D64080E450D2A286F1A3E3FF73F1F260F003F;
defparam sp_inst_1.INIT_RAM_2B = 256'hC0000E7717F3820DC7924E72FE017A9F07EACD3953800CA6FBC36300200BA00F;
defparam sp_inst_1.INIT_RAM_2C = 256'h00001441609E9A60F3BB393344C8687D8E35F30384000E62D00715408003E003;
defparam sp_inst_1.INIT_RAM_2D = 256'h000037B6EC6768393ED7F69985679CC0CAC2661EC00003FD8707C88B80012400;
defparam sp_inst_1.INIT_RAM_2E = 256'h000024D6D860FEA56DA51FACCD32ED38FC21ADC5C01D017CBF03CF47C400EF00;
defparam sp_inst_1.INIT_RAM_2F = 256'h000030DEB0EAAFC92C8B166C1F931B007F60BDD6017F60C6C9C9F90BC6007600;
defparam sp_inst_1.INIT_RAM_30 = 256'h000040A9D006806515E8AD29CF10E8BF35EEE4288F802F5F31777905DC000000;
defparam sp_inst_1.INIT_RAM_31 = 256'h00080377E00B64799FFFD2B2574120CADDC7E72A17008F1F2288DE9054200000;
defparam sp_inst_1.INIT_RAM_32 = 256'h000001E02075C0BD3E3474E0B31ABDE0BE8F203A2E47FF9E80987E44C42C0000;
defparam sp_inst_1.INIT_RAM_33 = 256'h00000003C8E6083D42DE5671FABB87D03E2FACBC18E9FEF090DE7E0EDF488000;
defparam sp_inst_1.INIT_RAM_34 = 256'h00000401003FFD9BFBFF0071E1F0CD87FBA238D861D64EC61A660E70DF000000;
defparam sp_inst_1.INIT_RAM_35 = 256'h00000001A2CAA9A16FE86FE3D1492DF90288B054D3698167745F7E4469728000;
defparam sp_inst_1.INIT_RAM_36 = 256'h000000021AE087F3FD3AD7E0A16A40D59FB9503B1D2E01E8A24AB76EA67C8000;
defparam sp_inst_1.INIT_RAM_37 = 256'h00000000240C1DEC7B38B0D1C0408CF7ABBE92F238A0183D0C08DF911E685100;
defparam sp_inst_1.INIT_RAM_38 = 256'h00000001901A06D21DD754A0FE248A34D4CE47F670D48C9B3F0BBF063FF07200;
defparam sp_inst_1.INIT_RAM_39 = 256'h010000019E4014832C3D0561FDFF7BD8FA0FB2E068A50EA8D4243F8418D20B00;
defparam sp_inst_1.INIT_RAM_3A = 256'h070000007F0017553F3E64E16F41694476A26F2DECEBCBECD7117F092D6F1780;
defparam sp_inst_1.INIT_RAM_3B = 256'h1F0000001AA3BD90DFEC5EE16621E083F98A1E69EE364BF078E13F030CC44AE0;
defparam sp_inst_1.INIT_RAM_3C = 256'h7F8000000170882EEC03CD20682C684F6FF1B80307BC57BC411C94004C89F4F8;
defparam sp_inst_1.INIT_RAM_3D = 256'hFF0000001F04E30FA27AF1533CA0E4F0B1FA806A0F7E6EFC962F040028019DFE;
defparam sp_inst_1.INIT_RAM_3E = 256'hFF0000000F875BEE210233089B069B0364AFFE2A0FAC6497B1DCD58026A893FF;
defparam sp_inst_1.INIT_RAM_3F = 256'hFF000000138288B7CE0B2BE109F383477ACF8A28E5FF0139F8228C83AA860DFF;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[30:0],sp_inst_2_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 1;
defparam sp_inst_2.BLK_SEL = 3'b000;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFDC7FFEFDFFF4340000005FE181BFFEFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF5EFFFFDF5DA025020407B4798BFFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFF77FEFBFF6D34901C3011F2E101FFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_03 = 256'hFCFFFFFFFFFFFFFFFFFFFFFFFFFDFFB5FFEEFE258015677CCA5FFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_04 = 256'hF0FFFFFFFFFFFFFFFFFFFFFFFFFFAFFF6FDFFF7DC0C5FE4CDC3FFFFFFFFFFF3F;
defparam sp_inst_2.INIT_RAM_05 = 256'hC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFBED9BE02EFD9E64AFFFFFFFFFFF0F;
defparam sp_inst_2.INIT_RAM_06 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFDFFFF3FDF3DFFB733DED1AC08FFFFFFFFFFF03;
defparam sp_inst_2.INIT_RAM_07 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBBFBABDB0407DFFFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_08 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFBFE6421817FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_09 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBFFCD83C96BFFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0A = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF7FFFFDDC081FFFFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0B = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFD71071EFFFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0C = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2DF3B037FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0D = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFF590EE067FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0E = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFA729D99F5FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_0F = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFE0E7E0877FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_10 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40B98E705FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_11 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7FFFB7F08F9E3FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_12 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF27A09EC33FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_13 = 256'h01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF27C07BF77FFFFFFFFFF00;
defparam sp_inst_2.INIT_RAM_14 = 256'h07FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4F829E047FFFFFFFFFF80;
defparam sp_inst_2.INIT_RAM_15 = 256'h1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB7C0E7F373FFFFFFFFFFE0;
defparam sp_inst_2.INIT_RAM_16 = 256'h7FFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFEFA124E67FFFFFFFFFFFF8;
defparam sp_inst_2.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4808113FFFFFFFFFFFE;
defparam sp_inst_2.INIT_RAM_18 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFEFC3E3D13BFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F1B8FF771FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCB6EF4FEF25FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1F3F8DF641FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB5FBA027291FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FC841E0481FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7E38007E5CEFFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDCE042FC103FFFFFFFFFEFF;
defparam sp_inst_2.INIT_RAM_20 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC8BB1C3E8862FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDEE731FFE81BFFFFFFFFFDFF;
defparam sp_inst_2.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8FF806FFFFE5FFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_23 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0CD3807FFE7EBFFFFFFFFFFF;
defparam sp_inst_2.INIT_RAM_24 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF2C5EA81F783EFFFFFFFFBFFF;
defparam sp_inst_2.INIT_RAM_25 = 256'hFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFED2ED888FF3FF9FFFFFFFBCFF;
defparam sp_inst_2.INIT_RAM_26 = 256'hF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC59E0C01FC62FFFFFFFFE53F;
defparam sp_inst_2.INIT_RAM_27 = 256'hC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9067DF81F5C01FFFFFFFFFF0F;
defparam sp_inst_2.INIT_RAM_28 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF84BFB83983F85FFFFFFFF7303;
defparam sp_inst_2.INIT_RAM_29 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF65DFF03803C6DFFFFFFFFFE00;
defparam sp_inst_2.INIT_RAM_2A = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF419FC20800E1BFFFFFFFFBE00;
defparam sp_inst_2.INIT_RAM_2B = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE413F0603F83267FFFFFBF7F00;
defparam sp_inst_2.INIT_RAM_2C = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC1763B9DB1FEEFFFFFFDFFE00;
defparam sp_inst_2.INIT_RAM_2D = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8E3F1DC00061E1BFFFF7FB8B00;
defparam sp_inst_2.INIT_RAM_2E = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9236BC80E1FF0F2FFFFFFDFF00;
defparam sp_inst_2.INIT_RAM_2F = 256'h00DDDCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB5C3FF80F077F824FFFFF77FE00;
defparam sp_inst_2.INIT_RAM_30 = 256'h0021FFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9B81DC00448E001FFF7FD7FFF00;
defparam sp_inst_2.INIT_RAM_31 = 256'h00FF31F3FFFFFFFFFFFFFFFFFFFFFFFFFFFFF19A1FC342E40003FFFFFF58FB00;
defparam sp_inst_2.INIT_RAM_32 = 256'h00B8610EFFFFFFFFFFFFFFFFFFFFFFFFF7FFF8F83F466FFC2042FFFFFFD6FE00;
defparam sp_inst_2.INIT_RAM_33 = 256'h0099FCFF7FFFFFFFFFFFFFFFFFFFFFFFFBFFFAE05E5CB7FE7FC37FFFFF2EDF00;
defparam sp_inst_2.INIT_RAM_34 = 256'h007FF37CDFFFFFFFFFFFFFFFFFFFFFFFFFFFA4C83FB8E7DC11FDFFFFFF7FD600;
defparam sp_inst_2.INIT_RAM_35 = 256'h0161B07FB7FFFFFFFFFFFFFFFFFFFFFFFFFFFD601F63018780241FFFFF87CB00;
defparam sp_inst_2.INIT_RAM_36 = 256'h07FB9FFE65FFFFFFFFFFFFFFFFFFFFFFFFFDF7000F0C00077FFC1FFFFFFEE980;
defparam sp_inst_2.INIT_RAM_37 = 256'h1FF41F999B7FFFFFFFFFFFFFFFFFFFFFFFFBEC060E884016FFFFFFFDF3EDFBE0;
defparam sp_inst_2.INIT_RAM_38 = 256'h7F1FF031F2EFFFFFFFFFFFFFFFFFFFFFFDF6BFC03C00008FC3F3FF7FBFFF7FF8;
defparam sp_inst_2.INIT_RAM_39 = 256'hFFFFC3FFFCB7FFFFFFFFFFFFFFFFFFFFFFE775207AA0081807F3FFFE797D7AFE;
defparam sp_inst_2.INIT_RAM_3A = 256'hFFFF1FFF92ECFFFFFFFFFFFFFFFFFFFFFB003CA0FE02719C07FFFFFFFECCF1FF;
defparam sp_inst_2.INIT_RAM_3B = 256'hFF7C1E7FFC7A3FFFFFFFFFFFFFFFFFFEFA001C02B612009E07F5FFFEDDFF83FF;
defparam sp_inst_2.INIT_RAM_3C = 256'hFFFABC7FFFEE0FFFFFFFFFFFFFFFF3E7F60010097E0B056E0FF3FFFFFFFC77FF;
defparam sp_inst_2.INIT_RAM_3D = 256'hFFF951F16FE3FBFFFFFFFFFFFFFBFFD79FA000005C8412FE0FF3FFFFFFF906FF;
defparam sp_inst_2.INIT_RAM_3E = 256'hFFB98E05EFFDD7FFFFFFFFFFFFFFB7B325BE0021140C00DC4FFBFFFFFEFCBDFF;
defparam sp_inst_2.INIT_RAM_3F = 256'hFFFE0BBF1A7DDD3FFFFFFFFF7FFFDA6B03ED00715CA1041CFE1CFFFFF79A1CFF;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[30:0],sp_inst_3_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 1;
defparam sp_inst_3.BLK_SEL = 3'b001;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'hFF740FF5FBFFFF1FFFFFFFF9FF7FF024001700000FFC4C19F80C7FFFFFF77CFF;
defparam sp_inst_3.INIT_RAM_01 = 256'hFFF81F03A3FFFF87FFFFEF917FB7F00A004E022286A00E6380042FFFFFEFAEFF;
defparam sp_inst_3.INIT_RAM_02 = 256'hFF181FC087FEDF10FFFFFF00FF37F075000108272E67395304063FFFFEF7F9FF;
defparam sp_inst_3.INIT_RAM_03 = 256'hFF3837900FE587D8FFFFFF907707F031000480173DCE78040C043FFFFABDEEFF;
defparam sp_inst_3.INIT_RAM_04 = 256'hFF3067818215FF051FDFFAFCBC01F8E20000A114BFAE6F0CD0013FEFFDB19DFF;
defparam sp_inst_3.INIT_RAM_05 = 256'hFF2463039063E3C3C7D768FCBC00D87C0020E01AAAC27B10A1001FFFE9F6A0FF;
defparam sp_inst_3.INIT_RAM_06 = 256'hFF04001A0B43C9DCB77F18FC5401F87C0003061AA00E4B9002012FFFFE567AFF;
defparam sp_inst_3.INIT_RAM_07 = 256'hFC38161594C45FCC59ED64F87607FC780001C755A08C9F1D00006FFFF38AF9FF;
defparam sp_inst_3.INIT_RAM_08 = 256'hF017269BE2101BE0EF761000371EFC7001087319737D298400083FFFFE66E73F;
defparam sp_inst_3.INIT_RAM_09 = 256'hC08F6FFF3408333507C8C080371478780421A3C91E6FC2C150B01FFEF9BDEF0F;
defparam sp_inst_3.INIT_RAM_0A = 256'h008F7EFF50FD87E127C500801F483C7C029758A578FF9C9E00B93FFFFA31CB03;
defparam sp_inst_3.INIT_RAM_0B = 256'h00CC0BFFC1C2DFFC02E202201E105C7E0032919B3ABDF84008695BFFEF4CFB00;
defparam sp_inst_3.INIT_RAM_0C = 256'h00C078D9FB11FFFF00F182E024DE2C7E0122AD13DC12F51334B21FFFFE7BD500;
defparam sp_inst_3.INIT_RAM_0D = 256'h00E24040A7C3F63F814D8FE1109F1631E3AA6DA26C866FA62247BFFFEF75ED00;
defparam sp_inst_3.INIT_RAM_0E = 256'h00F191853F0B07FF26071FE054FB5E1095A038D179DE4FEDDEA73FFF8DAA6200;
defparam sp_inst_3.INIT_RAM_0F = 256'h00FDC505FC800BFF920036404E121C47B6409819B8C83E1B1FF7FFFFFEDF7400;
defparam sp_inst_3.INIT_RAM_10 = 256'h00F8870FE16000FF408069405C0E1C4018980941268D15978181FFFFFB4EB300;
defparam sp_inst_3.INIT_RAM_11 = 256'h00F8EB8FC2C188FFA10098000C1EBC08FE583164759536AB03027FFFFDF36800;
defparam sp_inst_3.INIT_RAM_12 = 256'h00FEE107851F5FFFC002DA00041C781D902BC0724684A4BE5F007FFF7E97FF00;
defparam sp_inst_3.INIT_RAM_13 = 256'h00FC6B16043C0CDF3281840C0C18ED0EDC6E8D30683691D2FE55FFFFD47BFF00;
defparam sp_inst_3.INIT_RAM_14 = 256'h00FCF228186007FFEC81CC001E0B682E840AAFC19830173F3E4FFFFFF1DFFF00;
defparam sp_inst_3.INIT_RAM_15 = 256'h00FF945830D417FDF9B100001E0A06F3040C8CC042043F5F153FFBFFAD4AFF00;
defparam sp_inst_3.INIT_RAM_16 = 256'h00FE3198257C405FE520D0005D0116BDFE490C435A01AB480BD7FFFD340FF600;
defparam sp_inst_3.INIT_RAM_17 = 256'h01FFAFD9005B100F7030900078CF8FBAC7CC0C315C101A424ABFF7FFFF4EF600;
defparam sp_inst_3.INIT_RAM_18 = 256'h07FFA7C88266C30F9CB80000DA4B938382B8017C50001160B3BFBFFFFDAFFA80;
defparam sp_inst_3.INIT_RAM_19 = 256'h1FFFB780A8DD212FCD1800D367E2D31C043402B6A8000444DAAFBFFDFF6FFFE0;
defparam sp_inst_3.INIT_RAM_1A = 256'h7FFD8E08F1F00006E1A000C6213EB07E02B4459BC400050C7CEFFEF7FA5FFBF8;
defparam sp_inst_3.INIT_RAM_1B = 256'hFFFF6A0B64E10418764079B62338816200A4014FB0001D4A82BF9DCFFF23F9FE;
defparam sp_inst_3.INIT_RAM_1C = 256'hFFFF3003BB8E80107DC0A1BE61AA09780FAC01E64400250C0203FF2BDFCDF9FF;
defparam sp_inst_3.INIT_RAM_1D = 256'hFFFF2011770002A74DEB7B9D150B0C99097E017688018900AC8FF2FFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_1E = 256'hFFFEFC07730004DE7FD1CD39680F0D031D9C018EC001170E8C55FBEBFF7FFFFF;
defparam sp_inst_3.INIT_RAM_1F = 256'hFFFFE80EE202154F6473BD5DF2FC0904054B031E68018690329DE350FFFFFFFF;
defparam sp_inst_3.INIT_RAM_20 = 256'hFFFFD7CB8800325F0625919431030F220C1F005F800DDE9141188AF2FFFFFFFF;
defparam sp_inst_3.INIT_RAM_21 = 256'hFFFFFDCB30040E2F23E5730920DE0518022A8017290F5CC3E44190FFFFFFFFFF;
defparam sp_inst_3.INIT_RAM_22 = 256'hFFFFFC56571CA0F4DEBC7C8C903C41060A0FC02B643E620ED7C5C9F8FFFC6FFF;
defparam sp_inst_3.INIT_RAM_23 = 256'hFFFFFFB8AA7DA37FEEE3215D4065D29C03ADC032A8BE6D5CD5002BC0FF7003FF;
defparam sp_inst_3.INIT_RAM_24 = 256'hFFFFFD9064C2F11D3FF02D177A00E08602B5401013F7DCF06FA1B6A87F0003FF;
defparam sp_inst_3.INIT_RAM_25 = 256'hFFFFFDA0C384F0CD5A323F09DE0D28720B8940342B1D8C3040D5AD7C7F001BFF;
defparam sp_inst_3.INIT_RAM_26 = 256'hFFFFFA81CF87DFCBDF5A36624A0F8C722CD8606407562D1C86FD183C1FE83FFF;
defparam sp_inst_3.INIT_RAM_27 = 256'hFFFFFF9F3F80B64CFE5767815E07040E0896607C677966814F7B24641BF93FFF;
defparam sp_inst_3.INIT_RAM_28 = 256'hFFFFFF3ADFC163DB53F1B502320BB00E08F2A014BE2DE1620F0396181BF81FFF;
defparam sp_inst_3.INIT_RAM_29 = 256'hFCFFF9D3DB9751EF88089E893B0D501C0316980C4F3F6A183409C3C00FF808FF;
defparam sp_inst_3.INIT_RAM_2A = 256'hF0FFF9C7FFFE0D7F9BE8A681D108E81107C20801CB80E601DC00D61F27FF003F;
defparam sp_inst_3.INIT_RAM_2B = 256'hC0FFF64D6FFC57FBD8600401818CF43703150805100003E17C00E30027FFA00F;
defparam sp_inst_3.INIT_RAM_2C = 256'h00FFFC879F717995BC418A01FA06F3700C620408080001FDEC00F14083FFE003;
defparam sp_inst_3.INIT_RAM_2D = 256'h00FFFFB5104393E375284D00FA01211F8E0D840CD00000FDF800389803FFE400;
defparam sp_inst_3.INIT_RAM_2E = 256'h00FFFF482010F95633C694011A40B8FE41ACD43DE00000FF40003F0047FFEF00;
defparam sp_inst_3.INIT_RAM_2F = 256'h00FFFEB24010AF3E3B2DD9020C209CDEC9AE162EC0FF803EF000050847FFFF00;
defparam sp_inst_3.INIT_RAM_30 = 256'h00FFFF272002FC90FA186AC240A0176AB2B30B980380303FFC800701DCFFFF00;
defparam sp_inst_3.INIT_RAM_31 = 256'h00FFFEEF000B9F8FE0023441E9D01B76535481D90F0008F378600380F0FFFF00;
defparam sp_inst_3.INIT_RAM_32 = 256'h00FFFDDC4071F8BD41C279012B518E75A343A0FA1E400470F16801C40FFFFF00;
defparam sp_inst_3.INIT_RAM_33 = 256'h00FFFBBC00E0F10FBD20E980375291326037A8BC781A033F00C001C01F4FFF00;
defparam sp_inst_3.INIT_RAM_34 = 256'h00FFFFFC003FF06704014380E668A96900BE38DCE1ACB03FE24401801FCFFF00;
defparam sp_inst_3.INIT_RAM_35 = 256'h00FFFFFE22EAB8B690124201167FD127D17FB049C301FE078E0801C479F3FF00;
defparam sp_inst_3.INIT_RAM_36 = 256'h00FFFFFE3BE1761E02066A013E7D4D2EEC77F011030FFE15E82300E027F03F00;
defparam sp_inst_3.INIT_RAM_37 = 256'h00FFFFFC3FFFCF87849D09001CD0270F4C437032078FFFDDF1FB00700E607F00;
defparam sp_inst_3.INIT_RAM_38 = 256'h00FFFFFF9FE7A439E234BB400A944948C3E1E06207ABFFAF53E640FC1FF01F00;
defparam sp_inst_3.INIT_RAM_39 = 256'h01FFFFFF9FFFB0C7D3C0EB801A0CD1AF4FF271641F8AFFDCDA67C07C1FC02F00;
defparam sp_inst_3.INIT_RAM_3A = 256'h07FFFFFF1FFFA624C0C5AB00034FC13EFB5FE00413FC7F9CD3F780FF0B6F4780;
defparam sp_inst_3.INIT_RAM_3B = 256'h1FFFFFFF6FDE92AF3007D8006F7DFAD73E770140118C3F8C7BA2C0FF0BC44BE0;
defparam sp_inst_3.INIT_RAM_3C = 256'h7F7FFFFF8F7FF4F113FE47C0595D9E75972D8748F0003F8C0EFFEFFF07CFF0F8;
defparam sp_inst_3.INIT_RAM_3D = 256'hFFFFFFFFCCFCD9F07DF4746055DDFF6FDE469F09F8801ECC3B41E7FFEE5E7DFE;
defparam sp_inst_3.INIT_RAM_3E = 256'hFFFFFFFFF07E481B16EF4E313FF9815715F71F09F0001CE4377135FFE7EF73FF;
defparam sp_inst_3.INIT_RAM_3F = 256'hFFFFFFFFFC7D06C8ADFA1270FF4DDEBBCD766B8BFA0079C823FD7DFC657FFFFF;

SP sp_inst_4 (
    .DO({sp_inst_4_dout_w[30:0],sp_inst_4_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]})
);

defparam sp_inst_4.READ_MODE = 1'b0;
defparam sp_inst_4.WRITE_MODE = 2'b00;
defparam sp_inst_4.BIT_WIDTH = 1;
defparam sp_inst_4.BLK_SEL = 3'b000;
defparam sp_inst_4.RESET_MODE = "SYNC";
defparam sp_inst_4.INIT_RAM_00 = 256'hFF000000000000000000000023800102000BCBFFFFFFA07E7FC00100000000FF;
defparam sp_inst_4.INIT_RAM_01 = 256'hFF00000000000000000000000A1000020A25FDAFDFBF84F867C00000000000FF;
defparam sp_inst_4.INIT_RAM_02 = 256'hFF000000000000000000000008801040092CB6FE3CFEE171EFE00000000000FF;
defparam sp_inst_4.INIT_RAM_03 = 256'hFC00000000000000000000000002004A001101DA7FEA9BE335E00000000000FF;
defparam sp_inst_4.INIT_RAM_04 = 256'hF0000000000000000000000000005000902000823F3A07B3E3E000000000003F;
defparam sp_inst_4.INIT_RAM_05 = 256'hC0000000000000000000000000000000C00412641FD10E639B7000000000000F;
defparam sp_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000020000C020C20048CC21EE73F70000000000003;
defparam sp_inst_4.INIT_RAM_07 = 256'h000000000000000000000000000000000000004404543CFFF830000000000000;
defparam sp_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000004000000004039BDFFF8000000000000;
defparam sp_inst_4.INIT_RAM_09 = 256'h00000000000000000000000000000000000000002400727FF69C000000000000;
defparam sp_inst_4.INIT_RAM_0A = 256'h00000000000000000000000000000000000002080000E23F7E1C000000000000;
defparam sp_inst_4.INIT_RAM_0B = 256'h00000000000000000000000000000000000000002000E8EFFE1C000000000000;
defparam sp_inst_4.INIT_RAM_0C = 256'h00000000000000000000000000000000000000000001D20FFFCC000000000000;
defparam sp_inst_4.INIT_RAM_0D = 256'h00000000000000000000000000000000000008000003E6FFFF9C000000000000;
defparam sp_inst_4.INIT_RAM_0E = 256'h00000000000000000000000000000000000001400007CD7FE60E000000000000;
defparam sp_inst_4.INIT_RAM_0F = 256'h00000000000000000000000000000000000000040007F1FFFF8C000000000000;
defparam sp_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000FF07FF8FE000000000000;
defparam sp_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000048000CC0FFFE1C000000000000;
defparam sp_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000080001D85F7EFCC000000000000;
defparam sp_inst_4.INIT_RAM_13 = 256'h0100000000000000000000000000000000000000001D83FFBF8C000000000000;
defparam sp_inst_4.INIT_RAM_14 = 256'h0700000000000000000000000000000000000000003B07FFFFFC000000000080;
defparam sp_inst_4.INIT_RAM_15 = 256'h1F0000000000000000000000000000000000000000783FFFFF8C0000000000E0;
defparam sp_inst_4.INIT_RAM_16 = 256'h7F0000000000000000000000001000000000000000705FFFE7840000000000F8;
defparam sp_inst_4.INIT_RAM_17 = 256'hFF0000000000000000000000000000000000000000C03F7F81EC0000000000FE;
defparam sp_inst_4.INIT_RAM_18 = 256'hFF0000000000000000000000000000020000000000903C1FF1C40000000000FF;
defparam sp_inst_4.INIT_RAM_19 = 256'hFF000000000000000000000000000000000000000180E47FFF8E0000000000FF;
defparam sp_inst_4.INIT_RAM_1A = 256'hFF00000000000000000000000000000000000000030110BFEFDE0000000000FF;
defparam sp_inst_4.INIT_RAM_1B = 256'hFF000000000000000000000000000000000000000300C07FF7FE0000000000FF;
defparam sp_inst_4.INIT_RAM_1C = 256'hFF00000000000000000000000000000000000000040105FDF2EE0000000000FF;
defparam sp_inst_4.INIT_RAM_1D = 256'hFF000000000000000000000000000000000000000C037BFE04FE0000000000FF;
defparam sp_inst_4.INIT_RAM_1E = 256'hFF00000000000000000000000000000000000000181C7FFFE7FF0000000000FF;
defparam sp_inst_4.INIT_RAM_1F = 256'hFF000000000000000000000000000000000000001031FFFFC1FE0000000000FF;
defparam sp_inst_4.INIT_RAM_20 = 256'hFF000000000000000000000000000000000000003247E3FE887F0000000000FF;
defparam sp_inst_4.INIT_RAM_21 = 256'hFF000000000000000000000000000000000000002018CFFFE81E0000000000FF;
defparam sp_inst_4.INIT_RAM_22 = 256'hFF000000000000000000000000000000000000006007FFFFFFE50000000000FF;
defparam sp_inst_4.INIT_RAM_23 = 256'hFF00000000000000000000000000000000000000E02C7FFFFE7EC000000000FF;
defparam sp_inst_4.INIT_RAM_24 = 256'hFF00000000000000000000000000000000000000C0A11FFFF83F0000000000FF;
defparam sp_inst_4.INIT_RAM_25 = 256'hFC000000000000000000000000000000000000010912777FF3FE6000000000FF;
defparam sp_inst_4.INIT_RAM_26 = 256'hF0000000000000000000000000000000000000030261F3FFFFFF00000000003F;
defparam sp_inst_4.INIT_RAM_27 = 256'hC000000000000000000000000000000000000006000207FFFFFE00000000000F;
defparam sp_inst_4.INIT_RAM_28 = 256'h000000000000000000000000000000000000000600047FFFFFFA000000000003;
defparam sp_inst_4.INIT_RAM_29 = 256'h00000000000000000000000000000000000000080000FFFFFFF2000000000000;
defparam sp_inst_4.INIT_RAM_2A = 256'h00000000000000000000000000000000000000080203FFFFFFFE000000000000;
defparam sp_inst_4.INIT_RAM_2B = 256'h0000000000000000000000000000000000000018000FFFFF83FF800000000000;
defparam sp_inst_4.INIT_RAM_2C = 256'h0000000000000000000000000000000000000010009C0027000F000000000000;
defparam sp_inst_4.INIT_RAM_2D = 256'h000000000000000000000000000000000000003000E03FFFE001C00000000000;
defparam sp_inst_4.INIT_RAM_2E = 256'h000000000000000000000000000000000000002001437F1FFF00300000000000;
defparam sp_inst_4.INIT_RAM_2F = 256'h003DDF00000000000000000000000000000000200007F0FFFFFFF00000000000;
defparam sp_inst_4.INIT_RAM_30 = 256'h00E1FFE000000000000000000000000000000040023FFBB7FFFE000000000000;
defparam sp_inst_4.INIT_RAM_31 = 256'h00FFFFFC00000000000000000000000000000040003CBD1BFFFE000000000000;
defparam sp_inst_4.INIT_RAM_32 = 256'h00E79EFF0000000000000000000000000800010000B19003FFFF000000000000;
defparam sp_inst_4.INIT_RAM_33 = 256'h00E003078000000000000000000000000400010001A34801FFFE800000000000;
defparam sp_inst_4.INIT_RAM_34 = 256'h00800C83E000000000000000000000000000030000471823FFFE000000000000;
defparam sp_inst_4.INIT_RAM_35 = 256'h019FCF8078000000000000000000000000000200009CFE7FFFFFE00000000000;
defparam sp_inst_4.INIT_RAM_36 = 256'h07047C019E00000000000000000000000000080000F3FFFFFFFFE00000000080;
defparam sp_inst_4.INIT_RAM_37 = 256'h1F0FE066678000000000000000000000000002000177FFFFFFFC0000000000E0;
defparam sp_inst_4.INIT_RAM_38 = 256'h7FE00FCE01F0000000000000000000000000000003FFFF7FFFFC0000000000F8;
defparam sp_inst_4.INIT_RAM_39 = 256'hFF003C000078000000000000000000000000080005DFF7FFFFFC0000000000FE;
defparam sp_inst_4.INIT_RAM_3A = 256'hFF00E0007D1F000000000000000000000000000001FF8EFFFFF80000000000FF;
defparam sp_inst_4.INIT_RAM_3B = 256'hFF83E1800387C00000000000000000000000000009EFFFDFFFFA0000000000FF;
defparam sp_inst_4.INIT_RAM_3C = 256'hFF0743800001F00000000000000000180000000001FCFBFFFFFC0000000000FF;
defparam sp_inst_4.INIT_RAM_3D = 256'hFF06AE0E00003C00000000000000002C00400000037BEFFFFFFC0000000000FF;
defparam sp_inst_4.INIT_RAM_3E = 256'hFF467FFE10000E00000000000000004C004000002BF3FFFFFFFE0000000000FF;
defparam sp_inst_4.INIT_RAM_3F = 256'hFF01FBF0E58023C0000000000000001C004200002357FBFFFFFF0000000000FF;

SP sp_inst_5 (
    .DO({sp_inst_5_dout_w[30:0],sp_inst_5_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]})
);

defparam sp_inst_5.READ_MODE = 1'b0;
defparam sp_inst_5.WRITE_MODE = 2'b00;
defparam sp_inst_5.BIT_WIDTH = 1;
defparam sp_inst_5.BLK_SEL = 3'b001;
defparam sp_inst_5.RESET_MODE = "SYNC";
defparam sp_inst_5.INIT_RAM_00 = 256'hFF8BEFEA040000E0000000000000001E006000014003F3FFFFFF8000000000FF;
defparam sp_inst_5.INIT_RAM_01 = 256'hFF07FF7C7C000078000010000000001E00000001005FF3DFFFFFC000000000FF;
defparam sp_inst_5.INIT_RAM_02 = 256'hFFE7FFFFF80100AF000000000400000E000600008098C6AFFFFFC000000000FF;
defparam sp_inst_5.INIT_RAM_03 = 256'hFFC7F7EFF0180007800000000C00000E00032400003186FFFFFFC000000000FF;
defparam sp_inst_5.INIT_RAM_04 = 256'hFFCFAFFFFDEA0002E00000004000001C000100010001807BFFFEC000000000FF;
defparam sp_inst_5.INIT_RAM_05 = 256'hFFDBFFFFEF9C1C00380000004000000000010000000100EFFFFFE000000000FF;
defparam sp_inst_5.INIT_RAM_06 = 256'hFFFBFDFBFCBC36200C0000002800000000000000000180CFFFFFD000000000FF;
defparam sp_inst_5.INIT_RAM_07 = 256'hFCC7FFF7FBFBA00006000004080000000000000000030093FFFFF000000000FF;
defparam sp_inst_5.INIT_RAM_08 = 256'hF0E8FF9FFFEFE40000800000080000000020804400020023FFF7F0000000003F;
defparam sp_inst_5.INIT_RAM_09 = 256'hC070FFFF2BF7CC0000300000080004000018102400100406EF4FE0000000000F;
defparam sp_inst_5.INIT_RAM_0A = 256'h0070FFFFFF0EF80000380000201000000008120884000001FF46E00000000003;
defparam sp_inst_5.INIT_RAM_0B = 256'h00337BFFFE3DA000001C00002040000000850A44C4020003F796E00000000000;
defparam sp_inst_5.INIT_RAM_0C = 256'h003FFFD9FFEE0000000E00001000100000CD12E063680000CB4DE00000000000;
defparam sp_inst_5.INIT_RAM_0D = 256'h001DFF43FFFC0FC0000200002000080E1054925053718000DC98400000000000;
defparam sp_inst_5.INIT_RAM_0E = 256'h000E7F87FFF4F800000000002000001F685FC360D621A0002118400000000000;
defparam sp_inst_5.INIT_RAM_0F = 256'h000E3D07FFFFF400000008002008001C6CFF6361C33341E06000000000000000;
defparam sp_inst_5.INIT_RAM_10 = 256'h00077F0FFFFFFF00000000000010003FA667603A9130EE607E00000000000000;
defparam sp_inst_5.INIT_RAM_11 = 256'h00071F0FFFFE7700000060000000003F8027001A0200CD54FC00000000000000;
defparam sp_inst_5.INIT_RAM_12 = 256'h00031C07FFE0A000000020000000046FD804021802015B41A000000000000000;
defparam sp_inst_5.INIT_RAM_13 = 256'h00039017FFC3F320000000000000107D900162D806000E2D0000000000000000;
defparam sp_inst_5.INIT_RAM_14 = 256'h0003302FFF9FF8000000000000041473C0010030464008C0C000000000000000;
defparam sp_inst_5.INIT_RAM_15 = 256'h0001F05FFF3BE800000080000005107FE0000060A40000A0EA00040000000000;
defparam sp_inst_5.INIT_RAM_16 = 256'h0001F19FBEFFBFA0000000000286007A001000A0A4000435D600000000000000;
defparam sp_inst_5.INIT_RAM_17 = 256'h0100EFFF3FFCEFF0888000000780007D00100082200000199500080000000000;
defparam sp_inst_5.INIT_RAM_18 = 256'h0700BFFEFFFF3FF0600000002584007C01400083A80000030740000000000080;
defparam sp_inst_5.INIT_RAM_19 = 256'h1F00AFFCFEFEDFD0202400009C0400FA03C000431000000305C04000000000E0;
defparam sp_inst_5.INIT_RAM_1A = 256'h7F02BFF9FDFFFFF9101000001FC000F801C00044300000830BC00108000000F8;
defparam sp_inst_5.INIT_RAM_1B = 256'hFF00FFFBF8FEFBFF800000411FE000FC0BC00080480000017DC06230000000FE;
defparam sp_inst_5.INIT_RAM_1C = 256'hFF00FFF3B3F17FEF800010411FF000E60350000830000033F9FC00D4000000FF;
defparam sp_inst_5.INIT_RAM_1D = 256'hFF00DFF347FFFFD88000006049F0007E078800084000007F53780D00000000FF;
defparam sp_inst_5.INIT_RAM_1E = 256'hFF011FE713FFFFE00000024401F000FC07E80010100000F173BA0414000000FF;
defparam sp_inst_5.INIT_RAM_1F = 256'hFF001FEE23FDFAF018004220802204F80BF4000090026063CD7E1CBF000000FF;
defparam sp_inst_5.INIT_RAM_20 = 256'hFF002C0C07FFCFA000126201C0F000FC07F100006800000F9AFF750D000000FF;
defparam sp_inst_5.INIT_RAM_21 = 256'hFF0002680FFFFFD0D0128880D07102E405F50008D010A13C11BE6F00000000FF;
defparam sp_inst_5.INIT_RAM_22 = 256'hFF0003F21FFF7F0320408101E05902F007F50001B0001CF1003E3607000390FF;
defparam sp_inst_5.INIT_RAM_23 = 256'hFF0001F03FFFFF8000148C00B01A017206F60003500013EF2A7FD43F008FFCFF;
defparam sp_inst_5.INIT_RAM_24 = 256'hFF0003C07FFDFEE2000A0200903F007807FE0003E0002F1FF01FC95780FFFCFF;
defparam sp_inst_5.INIT_RAM_25 = 256'hFF0002C0FFFBFF00008D1002381F000C05FE8003C400F3FFF023D28380FFE4FF;
defparam sp_inst_5.INIT_RAM_26 = 256'hFF000501FFFFE00020871801AC1D400C03FF8003D821C7E37903E7C3E017C0FF;
defparam sp_inst_5.INIT_RAM_27 = 256'hFF00019FFF80C80031819800BE0EC02007FF80039880997FB004FB9BE406C0FF;
defparam sp_inst_5.INIT_RAM_28 = 256'hFF0003BFFFC1FC002C004800D704402007D7400340021E9DF04079E7E407E0FF;
defparam sp_inst_5.INIT_RAM_29 = 256'hFC00077FDFFFBE1037006000DF02A0220FF36003B00011E7C0003C3FF007F7FF;
defparam sp_inst_5.INIT_RAM_2A = 256'hF00006BFFFFFE000400010007F03102701BFF007F40001FFE00039E0D800FF3F;
defparam sp_inst_5.INIT_RAM_2B = 256'hC00009BF7FFFE804200838007F03000100EFF002EC00001F80001CFFD8005F0F;
defparam sp_inst_5.INIT_RAM_2C = 256'h00000373FFFFE40B000414003F81000301FFF807F800000000000EBF7C001F03;
defparam sp_inst_5.INIT_RAM_2D = 256'h0000005FFFBC0C0C801082003F80E02005FFF8032000000200000767FC001B00;
defparam sp_inst_5.INIT_RAM_2E = 256'h000000BFFFFF000FC0106100F780C00107DFF80200000000000000FFB8001000;
defparam sp_inst_5.INIT_RAM_2F = 256'h0000016DFFFF5007C01C2080F3C0E02100FFF80100000001060002F7B8000000;
defparam sp_inst_5.INIT_RAM_30 = 256'h000000D8FFFD0303000790003BC0A80148CCFC07007FC000020000FE23000000;
defparam sp_inst_5.INIT_RAM_31 = 256'h00000110FFF400C00007C9001BA0A401A4AA7E0600FFF00C8500007F0F000000;
defparam sp_inst_5.INIT_RAM_32 = 256'h00000223FF8E0742800184005DA0210240B85F0401BFF80F0E90003BF0000000;
defparam sp_inst_5.INIT_RAM_33 = 256'h00000443FF1F1FE00001D8004DA02A0981C8574007FBFC0FFF30003FE0B00000;
defparam sp_inst_5.INIT_RAM_34 = 256'h00000003FFC00F900000BC001F9336009041C7201E7EFF0FFDB8007FE0300000;
defparam sp_inst_5.INIT_RAM_35 = 256'h00000001DD154748000DF0006F902A0018004FB03CF9FF9FFBE6003B860C0000;
defparam sp_inst_5.INIT_RAM_36 = 256'h00000001C41E09E000C19C0057903A0010000FE0FCF1FF8DF79C001FD80FC000;
defparam sp_inst_5.INIT_RAM_37 = 256'h00000003C00030180063F60037B850A012000FC1F870FF85FE04000FF19F8000;
defparam sp_inst_5.INIT_RAM_38 = 256'h0000000060007BE4000BF00015F8168304101F81F8707FC77C1C0003E00FE000;
defparam sp_inst_5.INIT_RAM_39 = 256'h0100000060004F38001FF00005F00E0020000F83F0787FC4DF980003E03FF000;
defparam sp_inst_5.INIT_RAM_3A = 256'h07000000E00079F80003DC009CB0168100001FC3F00C3FC4D4080000F090F880;
defparam sp_inst_5.INIT_RAM_3B = 256'h1F000000F0016C400013D780988005288000FF87F0003FC4741F0000F03BB4E0;
defparam sp_inst_5.INIT_RAM_3C = 256'h7F000000708003C00001C6001680A18040027F87F0003FC418000000F8300FF8;
defparam sp_inst_5.INIT_RAM_3D = 256'hFF00000030030000000037800A00008000A17F87F0003E843090180011E002FE;
defparam sp_inst_5.INIT_RAM_3E = 256'hFF0000000001A404E810FFC0000066B88800FF87F8003C8C28060A0018100CFF;
defparam sp_inst_5.INIT_RAM_3F = 256'hFF0000000000F1067005FD80000020600081EB07F8003988440002001E0000FF;

SP sp_inst_6 (
    .DO({sp_inst_6_dout_w[30:0],sp_inst_6_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]})
);

defparam sp_inst_6.READ_MODE = 1'b0;
defparam sp_inst_6.WRITE_MODE = 2'b00;
defparam sp_inst_6.BIT_WIDTH = 1;
defparam sp_inst_6.BLK_SEL = 3'b000;
defparam sp_inst_6.RESET_MODE = "SYNC";
defparam sp_inst_6.INIT_RAM_00 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_01 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_02 = 256'hFF000000000000000000000000000000000000000000008000000000000000FF;
defparam sp_inst_6.INIT_RAM_03 = 256'hFC000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_04 = 256'hF00000000000000000000000000000000000000000000000000000000000003F;
defparam sp_inst_6.INIT_RAM_05 = 256'hC00000000000000000000000000000000000000000000000000000000000000F;
defparam sp_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000003;
defparam sp_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000001000000000000000;
defparam sp_inst_6.INIT_RAM_13 = 256'h0100000000000000000000000000000000000000000000004000000000000000;
defparam sp_inst_6.INIT_RAM_14 = 256'h0700000000000000000000000000000000000000000000000000000000000080;
defparam sp_inst_6.INIT_RAM_15 = 256'h1F000000000000000000000000000000000000000000000000000000000000E0;
defparam sp_inst_6.INIT_RAM_16 = 256'h7F000000000000000000000000000000000000000000000018000000000000F8;
defparam sp_inst_6.INIT_RAM_17 = 256'hFF00000000000000000000000000000000000000000000007E000000000000FE;
defparam sp_inst_6.INIT_RAM_18 = 256'hFF00000000000000000000000000000000000000000000000E000000000000FF;
defparam sp_inst_6.INIT_RAM_19 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_1A = 256'hFF000000000000000000000000000000000000000000000010000000000000FF;
defparam sp_inst_6.INIT_RAM_1B = 256'hFF000000000000000000000000000000000000000000000008000000000000FF;
defparam sp_inst_6.INIT_RAM_1C = 256'hFF00000000000000000000000000000000000000000000000D000000000000FF;
defparam sp_inst_6.INIT_RAM_1D = 256'hFF0000000000000000000000000000000000000000000001FB000000000000FF;
defparam sp_inst_6.INIT_RAM_1E = 256'hFF000000000000000000000000000000000000000000000018000000000000FF;
defparam sp_inst_6.INIT_RAM_1F = 256'hFF00000000000000000000000000000000000000000000003E000000000000FF;
defparam sp_inst_6.INIT_RAM_20 = 256'hFF000000000000000000000000000000000000000000000177800000000000FF;
defparam sp_inst_6.INIT_RAM_21 = 256'hFF000000000000000000000000000000000000000000000017E00000000000FF;
defparam sp_inst_6.INIT_RAM_22 = 256'hFF0000000000000000000000000000000000000000000000001A0000000000FF;
defparam sp_inst_6.INIT_RAM_23 = 256'hFF000000000000000000000000000000000000000000000001810000000000FF;
defparam sp_inst_6.INIT_RAM_24 = 256'hFF000000000000000000000000000000000000000000000007C00000000000FF;
defparam sp_inst_6.INIT_RAM_25 = 256'hFC00000000000000000000000000000000000000000000000C000000000000FF;
defparam sp_inst_6.INIT_RAM_26 = 256'hF00000000000000000000000000000000000000000000000000000000000003F;
defparam sp_inst_6.INIT_RAM_27 = 256'hC00000000000000000000000000000000000000000000000000000000000000F;
defparam sp_inst_6.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000003;
defparam sp_inst_6.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000007C00000000000000;
defparam sp_inst_6.INIT_RAM_2C = 256'h000000000000000000000000000000000000000000000000FFF0000000000000;
defparam sp_inst_6.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000001FFE000000000000;
defparam sp_inst_6.INIT_RAM_2E = 256'h00000000000000000000000000000000000000000000000000FFC00000000000;
defparam sp_inst_6.INIT_RAM_2F = 256'h0002200000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_30 = 256'h001E000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_35 = 256'h0100000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_6.INIT_RAM_36 = 256'h0700000000000000000000000000000000000000000000000000000000000080;
defparam sp_inst_6.INIT_RAM_37 = 256'h1F000000000000000000000000000000000000000000000000000000000000E0;
defparam sp_inst_6.INIT_RAM_38 = 256'h7F000000000000000000000000000000000000000000000000000000000000F8;
defparam sp_inst_6.INIT_RAM_39 = 256'hFF000000000000000000000000000000000000000000000000000000000000FE;
defparam sp_inst_6.INIT_RAM_3A = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_3B = 256'hFF000000000000000000000000000000000000000000002000000000000000FF;
defparam sp_inst_6.INIT_RAM_3C = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_3D = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_3E = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_6.INIT_RAM_3F = 256'hFF000400000000000000000000000000000000000000000000000000000000FF;

SP sp_inst_7 (
    .DO({sp_inst_7_dout_w[30:0],sp_inst_7_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]})
);

defparam sp_inst_7.READ_MODE = 1'b0;
defparam sp_inst_7.WRITE_MODE = 2'b00;
defparam sp_inst_7.BIT_WIDTH = 1;
defparam sp_inst_7.BLK_SEL = 3'b001;
defparam sp_inst_7.RESET_MODE = "SYNC";
defparam sp_inst_7.INIT_RAM_00 = 256'hFF001000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_01 = 256'hFF000080000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_02 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_03 = 256'hFF000800000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_04 = 256'hFF001000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_05 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_06 = 256'hFF000204000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_07 = 256'hFC000008000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_08 = 256'hF00000600000000000000000000000000000000000000000000000000000003F;
defparam sp_inst_7.INIT_RAM_09 = 256'hC0000000C000000000000000000000000000000000000000000000000000000F;
defparam sp_inst_7.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000003;
defparam sp_inst_7.INIT_RAM_0B = 256'h0000840000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0C = 256'h0000002600000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0D = 256'h000000BC00000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0E = 256'h0000007800000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_0F = 256'h000002F800000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_10 = 256'h000000F000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_11 = 256'h000000F000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_12 = 256'h000003F800000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_13 = 256'h000007E800000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_14 = 256'h00000FD000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_15 = 256'h00000FA000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_16 = 256'h00000E6040000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_17 = 256'h01001000C0000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_18 = 256'h0700400100000000000000000000000000000000000000000000000000000080;
defparam sp_inst_7.INIT_RAM_19 = 256'h1F004003010000000000000000000000000000000000000000000000000000E0;
defparam sp_inst_7.INIT_RAM_1A = 256'h7F004006020000000000000000000000000000000000000000000000000000F8;
defparam sp_inst_7.INIT_RAM_1B = 256'hFF000004070000000000000000000000000000000000000000000000000000FE;
defparam sp_inst_7.INIT_RAM_1C = 256'hFF00000C4C0000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_1D = 256'hFF00000CB80000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_1E = 256'hFF000018EC0000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_1F = 256'hFF000011DC0000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_20 = 256'hFF000033F80000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_21 = 256'hFF000017F00000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_22 = 256'hFF00000DE00000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_23 = 256'hFF00000FC00000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_24 = 256'hFF00003F800000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_25 = 256'hFF00003F000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_26 = 256'hFF00007E000000000000000010000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_27 = 256'hFF000060007F00000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_28 = 256'hFF000040003E00000000000008000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_29 = 256'hFC000000200000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_7.INIT_RAM_2A = 256'hF00000000000000000000000000000000000000000000000000000000000003F;
defparam sp_inst_7.INIT_RAM_2B = 256'hC00000008000000000000000000000000000000000000000000000000000000F;
defparam sp_inst_7.INIT_RAM_2C = 256'h0000000800000000000000000000000000000000000000000000000000000003;
defparam sp_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2E = 256'h0000000000000000000800000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000400000000000000000000;
defparam sp_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000F00000000000000000000;
defparam sp_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000600000000000000000000;
defparam sp_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000020000000000000000;
defparam sp_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000020000000000000000;
defparam sp_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000008000000000000000;
defparam sp_inst_7.INIT_RAM_39 = 256'h0100000000000000000000000000000000000000000000032000000000000000;
defparam sp_inst_7.INIT_RAM_3A = 256'h0700000000000000000000000000000000000000000800032800000000000080;
defparam sp_inst_7.INIT_RAM_3B = 256'h1F000000000000000000200000000000000000000000000380000000000000E0;
defparam sp_inst_7.INIT_RAM_3C = 256'h7F0000000000000000003800000000000000000000000003E0000000000000F8;
defparam sp_inst_7.INIT_RAM_3D = 256'hFF0000000000000000000800000000000000000000000103C0000000000000FE;
defparam sp_inst_7.INIT_RAM_3E = 256'hFF0000000000000000000000000000000000000000000303C0000000000000FF;
defparam sp_inst_7.INIT_RAM_3F = 256'hFF000000000000000000000000000000000014000000060780000000000000FF;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[30:0],sp_inst_8_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[0]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b00;
defparam sp_inst_8.BIT_WIDTH = 1;
defparam sp_inst_8.BLK_SEL = 3'b010;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'hFF00000001E2F9137EC80BF526990089628C0251C3FF9FF0FFFEC82206D851FF;
defparam sp_inst_8.INIT_RAM_01 = 256'hFF00000087650B4C6C3FE112D14ADCFFD59AE251F0731BEA3569EDF89F1C0BFF;
defparam sp_inst_8.INIT_RAM_02 = 256'hFF000000037554D5036FE4EA149EFBF9D1199357B069DFFB9DA0EF140A4A00FF;
defparam sp_inst_8.INIT_RAM_03 = 256'hFF00000001FBB7CE1C238023FB66590EBFE84C4B04FE2AE3A398E5C403CE01FF;
defparam sp_inst_8.INIT_RAM_04 = 256'hFF0000000119C54DDA600273C5CEBF2454BFBC8B05CD2287366E13B0800DE1FF;
defparam sp_inst_8.INIT_RAM_05 = 256'hFF000000008E46CED4430A04EAEBF48509F0B4AE00CA41AF7A6FA5FA88707BFF;
defparam sp_inst_8.INIT_RAM_06 = 256'hFF0000000119615B1A43307172762A697820BC0C2D78850FE92F7312B0CFD3FF;
defparam sp_inst_8.INIT_RAM_07 = 256'hFF200000006B5833B788C206814A465065F14E863863E61B38685DEC2B8FDEFF;
defparam sp_inst_8.INIT_RAM_08 = 256'hFF00000000150C035312F3E0B39192F2C5B8850E9BEC4EADC9CCF11F76EC70FF;
defparam sp_inst_8.INIT_RAM_09 = 256'hFF010000001ADCB1881506FC57F8F042D0EB874361D0694CA352B6238CF73FFF;
defparam sp_inst_8.INIT_RAM_0A = 256'hFF000000012D68080C2C13133DFE4052618C4EC3CE00978DC42807A09A80B6FF;
defparam sp_inst_8.INIT_RAM_0B = 256'hFC02000004AA9842385802219CA2B95AAE123981E7A46ECCA45F93B32A3B37FF;
defparam sp_inst_8.INIT_RAM_0C = 256'hF0420000103142893C427320EFC3BDCF90CFF11C136EF96B9238F57D19F4A93F;
defparam sp_inst_8.INIT_RAM_0D = 256'hC00000000BAC6CA61DB3418167410739D48B1102DFF80CC10EE1D37FB3D5F70F;
defparam sp_inst_8.INIT_RAM_0E = 256'h0000000004108E6FFC6FB9D3DB60095B05B3ED419EFF363D6EC810E7F3412A03;
defparam sp_inst_8.INIT_RAM_0F = 256'h000000005660112A8B9FBC5FEAB01B186702CC409C4092297201607E3B49BE00;
defparam sp_inst_8.INIT_RAM_10 = 256'h00000000BEA301FC899FBC95FD51CC486483D3820C6C6A6C3F30744281F87F00;
defparam sp_inst_8.INIT_RAM_11 = 256'h0000000068A53D801DFAFEB7F553ACEEE22D4BA065B2A864A6CB151C6FBD4E00;
defparam sp_inst_8.INIT_RAM_12 = 256'h0006002030028F081DC3DF75F97BA16FFC15B1F99FFAA1486E5B151636341C00;
defparam sp_inst_8.INIT_RAM_13 = 256'h00A01000C002C45C26435F7AFA23B7C3E86DD8F9EFF557D92637E3F6373B9600;
defparam sp_inst_8.INIT_RAM_14 = 256'h00040800768EF148ECE3FFBD7E3B00DD04F2C00D1F7A931DC36EFE91F4124500;
defparam sp_inst_8.INIT_RAM_15 = 256'h0045AA010399A3B577D38D7C7F3A0EC957FB2C07228D1EF57C88771D95180B00;
defparam sp_inst_8.INIT_RAM_16 = 256'h001AC20003476FFF47F3CEF27D308D784A33DA01EF146B873FABF904C035B800;
defparam sp_inst_8.INIT_RAM_17 = 256'h0016E00004007FA28EA1D2F07936300DE9DB4B87ADED71E2A7C4FF002064D000;
defparam sp_inst_8.INIT_RAM_18 = 256'h00854C005B03BDF5CFC4A7F4F93F36BF3387ABC7E88BD43A0998BFE024A0FE00;
defparam sp_inst_8.INIT_RAM_19 = 256'h00D020C0170099F98F206FF4FC39F86F4F032F878591E15D4308FFFF0E060E00;
defparam sp_inst_8.INIT_RAM_1A = 256'h001D2E240584F30D1BA07320F237F81D845D21F5E21D550F5EC37FE4DCDF1700;
defparam sp_inst_8.INIT_RAM_1B = 256'h01058240050159E28A0E0319F8DD97BCA0EED1A7F2B7884C66413FA7ECE47900;
defparam sp_inst_8.INIT_RAM_1C = 256'h0761DCA01F127DF13DF20CCBE4BE95E9EB88629DE156D90CA200FCD6FB47AB80;
defparam sp_inst_8.INIT_RAM_1D = 256'h1F1882900125180DDCDD0E05EFBC1285E6213F7565F2C56EB4793040EF02BAE0;
defparam sp_inst_8.INIT_RAM_1E = 256'h7FC8F9FE2001FF31BD8E80F0977F13113444BF77EE8CAD1527E3F385820C60F8;
defparam sp_inst_8.INIT_RAM_1F = 256'hFF01A57C2AE177EA5C9670074AF8130A480366F7D9CFF6B86B25B3525F8A45FE;
defparam sp_inst_8.INIT_RAM_20 = 256'hFF353DDA130133698709D8121CD809B6A463C37AFC567E6F4227F713FFCEEFFF;
defparam sp_inst_8.INIT_RAM_21 = 256'hFF524AE2B807E297DFC7EE143B892FB742AFE1EB36DAA2862C18E1C53FFE17FF;
defparam sp_inst_8.INIT_RAM_22 = 256'hFFF0BED407087793F199F8A378D9FF8FBB3B45FBC4048B13EE12BC248D741CFF;
defparam sp_inst_8.INIT_RAM_23 = 256'hFF077FF84F80FAF631867E9601FF5FB8516DA9E2591FCA2F700D8DC287731DFF;
defparam sp_inst_8.INIT_RAM_24 = 256'hFFAD7F5C578072DC086644AEDE7FF05122C3A0598EE5FACCC9EFF066D3C975FF;
defparam sp_inst_8.INIT_RAM_25 = 256'hFFDFEFFD4F8960DA61914171F13F3A120FA51006E0D617DB619B763E47C5FFFF;
defparam sp_inst_8.INIT_RAM_26 = 256'hFFFF5EA78485F294AF860182A4DFBB50408BF81443AF519467A06C776524BBFF;
defparam sp_inst_8.INIT_RAM_27 = 256'hFFEFFF7FE393F5AE929FF9DB043F6813B8FFC57F4332406925B8BFE86CC9FFFF;
defparam sp_inst_8.INIT_RAM_28 = 256'hFF5D7D5F8BE1FB9282BCE6D2E33FF41A1447A4EC3942287A48C10663134512FF;
defparam sp_inst_8.INIT_RAM_29 = 256'hFFEFBFFEF153FC287AE7C3A7CF3F40FAB8FFC360C9150B9FE003FE45121BC9FF;
defparam sp_inst_8.INIT_RAM_2A = 256'hFF5DB6A5B853F800FB9C0D8E887FECE4B070E2E9116197480FAFD9F30891A0FF;
defparam sp_inst_8.INIT_RAM_2B = 256'hFFEFDF95C05FFF45FF012D4D387D3728101146CF88C17FE5FE46A1789694BAFF;
defparam sp_inst_8.INIT_RAM_2C = 256'hFFFDCF7EE30FFDC7AF3D028B9216EC2FDD04850EC3A0166D86DDC897B33BBDFF;
defparam sp_inst_8.INIT_RAM_2D = 256'hFCDFFFFFEFCFF3E5E05DE95C222F3C21F6177C5B1142C3745FF9FD16B75380FF;
defparam sp_inst_8.INIT_RAM_2E = 256'hF0F7FFFECC3FFEFFC9E5C47C0DCFBA70119DFFC086003B69DF101637FD50813F;
defparam sp_inst_8.INIT_RAM_2F = 256'hC0FFFFFFB89FFFFF39E850957F3E9D462236A36406014706E701065E7517AD0F;
defparam sp_inst_8.INIT_RAM_30 = 256'h00FFFFFFBC2BDFFFF3C2D42569B86612923D61A24CE12968FEBAE1A83F70CE03;
defparam sp_inst_8.INIT_RAM_31 = 256'h00FFFFFFFE3B3FBFFC5E5D862402CD1AECEC38AFF3184CB81E90CE8DB3E85100;
defparam sp_inst_8.INIT_RAM_32 = 256'h00FFFFFFDF3F83C8EC6F846FB00726053F7C1C85C2F1C66D0E1CEE85F3852B00;
defparam sp_inst_8.INIT_RAM_33 = 256'h00FFFFFFDF33EBE7BF7EA0FBEF1E6303E60A001531DDDFE3BCC44378B1745B00;
defparam sp_inst_8.INIT_RAM_34 = 256'h00FFFFFFF9F7A38267C7BF9C7110A4C7B02203E501E2CBEB7B613B33C2267B00;
defparam sp_inst_8.INIT_RAM_35 = 256'h00FDFFFFEF86029F4A8C52F2BD172C076060594D2E63D9D8E83180F19C338E00;
defparam sp_inst_8.INIT_RAM_36 = 256'h00FFFFFFFB2308E7A805EBDCB4585E07706094F0B61BDD8706F82828B9DF0F00;
defparam sp_inst_8.INIT_RAM_37 = 256'h00FFFFEFF1A285EFF01F069228149E4B7C409B6F1BECB93299CD7FC3E28D4C00;
defparam sp_inst_8.INIT_RAM_38 = 256'h00FFFFFFFD8BB3A8E7AEC84FE58DA5930304F182D5F565AC55F4BF1AEBBD4700;
defparam sp_inst_8.INIT_RAM_39 = 256'h00FFFFFFBFD3F8F81C7C37C9FDDEB542828F68CEBECA3B5DE8F8631D707BDB00;
defparam sp_inst_8.INIT_RAM_3A = 256'h00DFFFFFFF917071CDF7329412FC7694D8EB2E29F1EB04572D03CC90FF862600;
defparam sp_inst_8.INIT_RAM_3B = 256'h00FFFFFFEF58704EC17F934E00192BCD2865E36E03E8C0065193918F2316F300;
defparam sp_inst_8.INIT_RAM_3C = 256'h00FFFFE7FC8321FD83E9E11A35A04139CE422CE4975D4E4D98EF709B02E35F00;
defparam sp_inst_8.INIT_RAM_3D = 256'h01FFFFFFBFC24003506FB7C2473A594F6BBBFC98F55F2BBDAE107F567604BF00;
defparam sp_inst_8.INIT_RAM_3E = 256'h07FFFFFFEDA7EC0B4A6F682926A0F17FA9F9DDF7E149FC23C37E594405937980;
defparam sp_inst_8.INIT_RAM_3F = 256'h1FFFFFFFBFE1F0A3D72C707F07A0221ED719DFDF83F4B6BE858924C9AE49E6E0;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[30:0],sp_inst_9_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b00;
defparam sp_inst_9.BIT_WIDTH = 1;
defparam sp_inst_9.BLK_SEL = 3'b010;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'hFFFFFFFFFE1CBEF2FF280FFAFF6FA6D4151CC3ABDC003F089CC139FDE35BDCFF;
defparam sp_inst_9.INIT_RAM_01 = 256'hFFFFFFFF789A7C4F8A4013FD78B5B6EE3C39E3A3DC007B991A8619FF71DFFBFF;
defparam sp_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFC8DB715187803F5DD6195F52FDD8225BF003F90260E1F1FFBEBFEFF;
defparam sp_inst_9.INIT_RAM_03 = 256'hFFFFFFFFFE09F131E0C4007FFBD9B7F6CB6E013507006B10BC47178FFFBFFFFF;
defparam sp_inst_9.INIT_RAM_04 = 256'hFFFFFFFFFEE5C3C18FF0000FC5F174C9E7BF01320621E300C193F3FF7FFDFDFF;
defparam sp_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFFD073744800003EAF57DEEE7E049108309C222C7EFE7FF7FF1FBFF;
defparam sp_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFEEBE22FFF800F80F079F10F80724191018784C9D7BE7713CFDBF5FF;
defparam sp_inst_9.INIT_RAM_07 = 256'hFFDFFFFFFFF917DE5C003FF8600DFC790296B308A07F0998C93E1FE037FFFCFF;
defparam sp_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFF77B260C01F3FF10036CF674BA7890400191BEB36CD718F6E678FF;
defparam sp_inst_9.INIT_RAM_09 = 256'hFFFEFFFFFFF33C0C400306FF8C01ABFF4C397A802E2FC766FA75B6200CC3FFFF;
defparam sp_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFDECE6790040313C400BFCD9E56318019FE0FFA3ED7379F057EBEFF;
defparam sp_inst_9.INIT_RAM_0B = 256'hFCFDFFFFFFDE34BC80080E21E05C5FA2522041E00DC83FB6FEA3F38C380C45FF;
defparam sp_inst_9.INIT_RAM_0C = 256'hF0BDFFFFEFDDB87040900F30F13CD3BD1D9080600081BC5073C79103E1F0AF3F;
defparam sp_inst_9.INIT_RAM_0D = 256'hC0FFFFFFFA507245E0103F98383E7EAFD77C9EFD0005F1E3F8BFF3007DC07F0F;
defparam sp_inst_9.INIT_RAM_0E = 256'h00FFFFFFFFE49477C1A0079C1C9FFC26F2FC17BF61E0CFFFB2FCC01800403B03;
defparam sp_inst_9.INIT_RAM_0F = 256'h00FFFFFFDF80139FF14043000C0FBE5C08FDC7AE001F2BBB9FFDE00401C61F00;
defparam sp_inst_9.INIT_RAM_10 = 256'h00FFFFFFFF739FD1F36043FA064F9C4F237CE46EEFFEFE82A1D47581FDF79800;
defparam sp_inst_9.INIT_RAM_11 = 256'h00FFFFFFEF727BCBF3650118060FD81C17FE647EE5FD419BDE7C1C8019B69C00;
defparam sp_inst_9.INIT_RAM_12 = 256'h00F9FFDFFFE0B0FFD37C00000227C1144AEF600740184577A0A0CCE9C7939C00;
defparam sp_inst_9.INIT_RAM_13 = 256'h005FEFFFFFE2EBE389FC0080030FC41285962006A02BDDCEE6107801D8F81600;
defparam sp_inst_9.INIT_RAM_14 = 256'h00FBF7FFFFF0FFB7815C40000317E02D5B0D100290957EFF0A6DAE9009F78C00;
defparam sp_inst_9.INIT_RAM_15 = 256'h00BA55FFFFF5FC03084C00020217EC0918823800D2B248FB837BCFFC07FB8F00;
defparam sp_inst_9.INIT_RAM_16 = 256'h00E53DFFFFF89003384C000202036E08F5C41C002031A9FE4058477CC7F04800;
defparam sp_inst_9.INIT_RAM_17 = 256'h00E91FFFFFF8401E785E0000020C7B014E243C00402B6FF1543380FFEFF31F00;
defparam sp_inst_9.INIT_RAM_18 = 256'h007AB3FFDFFFC014341B0000020758B904686C000CF7ECEDE50F401FFB871F00;
defparam sp_inst_9.INIT_RAM_19 = 256'h002FDF3FF7FCA038743F88040607D86003FCED0065EF78F3B5BE8000F1860F00;
defparam sp_inst_9.INIT_RAM_1A = 256'h00E2D1DBFFFC80F2FE0F8008040008003EA22F001E1093189E7D801B23CF1F00;
defparam sp_inst_9.INIT_RAM_1B = 256'h01FA7DBFFFFC60F87D97E3080C000F821F111E401CE16BF31A32C05812047F00;
defparam sp_inst_9.INIT_RAM_1C = 256'h079E235FFFFCC1F03E07F0C808000DC017F47C60333593F755FF03F907044380;
defparam sp_inst_9.INIT_RAM_1D = 256'h1FE77D6FFFFDE2CF3DA7F00210000F811BFC38081F7977310386FFFF1F01BFE0;
defparam sp_inst_9.INIT_RAM_1E = 256'h7F370601DFFD82E3FD73FF0F20800F20CFF83C0C1187574A001FFF1E7F8BAFF8;
defparam sp_inst_9.INIT_RAM_1F = 256'hFFFE5A83DBFF80F4FCA9FFF807800B483FFC3C0907813E4F90DFF073A70A07FE;
defparam sp_inst_9.INIT_RAM_20 = 256'hFFCAC225F3FFC1EE3F564FFD0CA01D715BDC5E8607CA09C5B7DFE013FFDE0EFF;
defparam sp_inst_9.INIT_RAM_21 = 256'hFFADB51D5FF985EA3FF817E058F01FB0FDD07E144F993A0C2FF8E0053FFE17FF;
defparam sp_inst_9.INIT_RAM_22 = 256'hFF0F412BFFF780FC03FA000067A00F8C65D41A067B27F7406FF283C0007C1FFF;
defparam sp_inst_9.INIT_RAM_23 = 256'hFFF88007BFFF0169458C80021E802FF8AF967E068F70E6401FFC622387F321FF;
defparam sp_inst_9.INIT_RAM_24 = 256'hFF5280A3BFFF83637667A2C03E800FD0DD3C2FA506B60F207E6000F6FFC687FF;
defparam sp_inst_9.INIT_RAM_25 = 256'hFF201002BFF78066E0EFFF9FF3C007F1F25A1FFE849E08037F84020187C23FFF;
defparam sp_inst_9.INIT_RAM_26 = 256'hFF00A1587CFA01FB7079DE7E842007F3BB742FEC8F6CCBB87FA0138847233BFF;
defparam sp_inst_9.INIT_RAM_27 = 256'hFF1000801FFC01DBE6F2002702C087F0470047FF8EE3C00A3F80000C2FC7BFFF;
defparam sp_inst_9.INIT_RAM_28 = 256'hFFA282A07FFE00FB1B8F3DF67DC003F9EBB027EC60BC1879F800FF8013421EFF;
defparam sp_inst_9.INIT_RAM_29 = 256'hFF1040010FFC00F786ECCFBD85C08718070007E032FA803FE00001BA3200DCFF;
defparam sp_inst_9.INIT_RAM_2A = 256'hFFA2495A47EC00FF04EB5BB390C003180F8F03F82EBE64080FA02601F80B9FFF;
defparam sp_inst_9.INIT_RAM_2B = 256'hFF10206A3FF000BA00DFFF75B601C0D86FEA878C573EC045FFC15E7B703C78FF;
defparam sp_inst_9.INIT_RAM_2C = 256'hFF0230811FF0007850E0FFB7CDE993DC23F807C23F7F060207C1FF979BE472FF;
defparam sp_inst_9.INIT_RAM_2D = 256'hFC20000013F0001A7FA0EB5705D1C3D8099773D6FFEFD5500FFEFC9E74DC3FFF;
defparam sp_inst_9.INIT_RAM_2E = 256'hF008000133C001003F15F924F7B1C1880E7D0055FF3F12F9FC1FF625FB60FF3F;
defparam sp_inst_9.INIT_RAM_2F = 256'hC000000047E00000FA1FE87EF7C022BC2DFD7CE3FFA1B0FFFFFFC42000E03D0F;
defparam sp_inst_9.INIT_RAM_30 = 256'h0000000043C020000F98B7B4750679EDE3F37E41C7E5E51E80397E0FEF3F7103;
defparam sp_inst_9.INIT_RAM_31 = 256'h0000000001C0C0401E2C97B55BFE73EEFF1C3F13F3A6DC80DBD87FC9BDC87000;
defparam sp_inst_9.INIT_RAM_32 = 256'h0000000020C07C371110C5E947F759FFC0FC1F70C50F8011901B4107FC703800;
defparam sp_inst_9.INIT_RAM_33 = 256'h0000000020CC141840F9CAE9F7EC7FFC1A0C0FB1026A4003A1469C878F834400;
defparam sp_inst_9.INIT_RAM_34 = 256'h0000000006087C7DB8393D26EFFC7BF8700220F8E1A5F86AA87E3DCF8FFE7800;
defparam sp_inst_9.INIT_RAM_35 = 256'h000200001079FD60B5DB1F31F9F07FF8E00006B0C27066CC0FC1FF0F7FFC0000;
defparam sp_inst_9.INIT_RAM_36 = 256'h0000000004DFF71857A89E4425F07FF8F0008EDF481BDF27F8FFD7D67FE7FC00;
defparam sp_inst_9.INIT_RAM_37 = 256'h000000100E5FFE100FFA959CACD01930FC0002C79BE571EEFE1680BC1E05FD00;
defparam sp_inst_9.INIT_RAM_38 = 256'h00000000027BFC571B8975AE1FC53F00FF1C8C7DD01C006FC64C801D343EFE00;
defparam sp_inst_9.INIT_RAM_39 = 256'h00000000402FFF07E78385D173D895810197543FEA58F741F03A9F834BFB3F00;
defparam sp_inst_9.INIT_RAM_3A = 256'h00200000000EFF8FF3002DFADFBC66A800F7191A7D0F1C248FFC3F800079D900;
defparam sp_inst_9.INIT_RAM_3B = 256'h0000000010BFFFB3FE806EF13F193896F0F3D816107AB006D2D8700023070000;
defparam sp_inst_9.INIT_RAM_3C = 256'h00000018037CFE0B9E101E69B9E840B600F1DB03E2B30E73E099F00C031FA000;
defparam sp_inst_9.INIT_RAM_3D = 256'h01000000443DBFFCF1D041EF9F380244C4401BE0147C2C63F06FFC2EF5FFC000;
defparam sp_inst_9.INIT_RAM_3E = 256'h07000000125C0FFCBF70C7FE1E70A2F3D2000A0E1801DFEFCC8BC8B807BC8080;
defparam sp_inst_9.INIT_RAM_3F = 256'h1F000000401E0FDC0E330E38BFA0B5D6590017207C070E5F05FF60E1D1EE99E0;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[30:0],sp_inst_10_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[2]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b00;
defparam sp_inst_10.BIT_WIDTH = 1;
defparam sp_inst_10.BLK_SEL = 3'b010;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'hFF0000000003400C00F7F000000018622863C307EC007F88C00006001C2423FF;
defparam sp_inst_10.INIT_RAM_01 = 256'hFF000000000183B071800C00060008100247E307DE007B09200006000E2004FF;
defparam sp_inst_10.INIT_RAM_02 = 256'hFF000000000208EAE78000002200000200238303BF007F00400000E0041401FF;
defparam sp_inst_10.INIT_RAM_03 = 256'hFF00000000060EFE0F38000004000001641201030780EB1040000870000000FF;
defparam sp_inst_10.INIT_RAM_04 = 256'hFF00000000023CBE300000003A0002160043010107C0E22100000C00000202FF;
defparam sp_inst_10.INIT_RAM_05 = 256'hFF0000000003F818BB00000015000210100C010183F7C06000101800000E04FF;
defparam sp_inst_10.INIT_RAM_06 = 256'hFF00000000061DF0040000000F8004B0178E010081FF804C004188EC003C08FF;
defparam sp_inst_10.INIT_RAM_07 = 256'hFF0000000006EFE1B00000001FF001AED16E0300607F009006C1E01FC00003FF;
defparam sp_inst_10.INIT_RAM_08 = 256'hFF000000000887DBF0000C000FFC01098B460100200001B00C9328E7091F87FF;
defparam sp_inst_10.INIT_RAM_09 = 256'hFF000000000C03E7B000F90003FE0400A3C7030010004379058A49DFF33C00FF;
defparam sp_inst_10.INIT_RAM_0A = 256'hFF0000000001F1986003FCEC03FF0022C1EA010004000FC00100C87FFFFF41FF;
defparam sp_inst_10.INIT_RAM_0B = 256'hFC0000000001E361C007F1DE03FF000DE1FE010003041F0101000C7FC7FFFAFF;
defparam sp_inst_10.INIT_RAM_0C = 256'hF00000000002079F800FE0CF00FF0000E3FF818000007E8F0C000EFFFE0F503F;
defparam sp_inst_10.INIT_RAM_0D = 256'hC0000000040F81FA000FC067C0FF81402BFF9F000003FE1C01000CFFFE3F800F;
defparam sp_inst_10.INIT_RAM_0E = 256'h00000000001F6398001FC063E07F83C8DDFFFA00001FF00011033FFFFFBFC403;
defparam sp_inst_10.INIT_RAM_0F = 256'h00000000201FEC60003F80F3F07FC1A3F7FF3811FFFFC44460021FFFFE3FE000;
defparam sp_inst_10.INIT_RAM_10 = 256'h00000000000C6002003F8011F83FE3B1DFFF0811EFFF1111420F8BFFFE0FE700;
defparam sp_inst_10.INIT_RAM_11 = 256'h00000000100F8004003F8001F83FE7E3E9FF8001E5FC762419BFE3FFFE4FE300;
defparam sp_inst_10.INIT_RAM_12 = 256'h00000000001F4000203F8001FC1FFEEBB77F8000C01F1ABC7FFFF3FFF86FE300;
defparam sp_inst_10.INIT_RAM_13 = 256'h00000000001D0000703F8001FC1FFBED7FFFC0006034203019EF87FFE007E900;
defparam sp_inst_10.INIT_RAM_14 = 256'h00000000000F0000703F8001FC0FFFF2FFFFE00070E001003D93C16FFE0FF300;
defparam sp_inst_10.INIT_RAM_15 = 256'h00000000000E0000F03FC001FC0FF3F6FFFDC00032C0B70000078003F807F000;
defparam sp_inst_10.INIT_RAM_16 = 256'h0000000000070000F03FE001FC0FF3F70FFFE0001FCF160000078083380FF700;
defparam sp_inst_10.INIT_RAM_17 = 256'h0000000000078001F03FC003FC03C7FEBFFFC0001FD0900C080F0000100FE000;
defparam sp_inst_10.INIT_RAM_18 = 256'h000000002000000BF83FF003FC00C746FFFFD0001300031012FF8000007FE000;
defparam sp_inst_10.INIT_RAM_19 = 256'h0000000008034007F81FF003F800079FFFFF90001A1086000E7F00000079F000;
defparam sp_inst_10.INIT_RAM_1A = 256'h000000000003000FFC1FFC07F80007FFFFFFD00001E22CE061FE00000030E000;
defparam sp_inst_10.INIT_RAM_1B = 256'h0100000000038007FE0FFC07F000007FFFFFE000010C940081FC000001FB8000;
defparam sp_inst_10.INIT_RAM_1C = 256'h070000000003020F3F0FFF37F000023FFFFF80000CE82C000800000000FBFC80;
defparam sp_inst_10.INIT_RAM_1D = 256'h1F00000000020133FD03FFFFE000007EFFFFC000008798C00000000000FFC0E0;
defparam sp_inst_10.INIT_RAM_1E = 256'h7F0000000002001FFD81FFFFC00000DFFFFFC000007828B0000000E00077D0F8;
defparam sp_inst_10.INIT_RAM_1F = 256'hFF0000000400000FFCC0FFFF800004B7FFFFC000007EC10400000F8C00F5F8FE;
defparam sp_inst_10.INIT_RAM_20 = 256'hFF0000000C000011FF603FFE0300020FFFFFA001003DFE3848001FEC0021F0FF;
defparam sp_inst_10.INIT_RAM_21 = 256'hFF00000000000005FFF00FF80700004FFFFF80038067DDF3D0071FFAC001E8FF;
defparam sp_inst_10.INIT_RAM_22 = 256'hFF00000000000000FFFC00009F000073FFFFE00180FB0CFF900D7FFFFF83E0FF;
defparam sp_inst_10.INIT_RAM_23 = 256'hFF00000000000000ED8F0001FF000007FFFFC001F08F11BFE003FFFC780CFEFF;
defparam sp_inst_10.INIT_RAM_24 = 256'hFF0000000000000081E7FD3FFF00002FFFFFD002F90FFC1F801FFF09E03FF8FF;
defparam sp_inst_10.INIT_RAM_25 = 256'hFF000000000000811F7FFFFFF200000FFFFFE0017F61FFFC807FFDFFF83FC0FF;
defparam sp_inst_10.INIT_RAM_26 = 256'hFF000000030000000C3FDFFE8700000FFFFFD003FFD3BC7F805FFFFFB8DFC4FF;
defparam sp_inst_10.INIT_RAM_27 = 256'hFF00000000000000190DFFFF0700000FFFFFB800FFFC3FF7C07FFFF3903FC0FF;
defparam sp_inst_10.INIT_RAM_28 = 256'hFF000000000000046473DB0DFE000007FFFFD813FFFFF78787FFFFFFECBFE1FF;
defparam sp_inst_10.INIT_RAM_29 = 256'hFF000000000000000113B0437A000007FFFFF81FFFFFFFC01FFFFFFFCDFF32FF;
defparam sp_inst_10.INIT_RAM_2A = 256'hFF000000000000000004E44C6F000007FFFFFC07FFFFFBF7F05FFFFE07F820FF;
defparam sp_inst_10.INIT_RAM_2B = 256'hFF000000000000000320038A4B800007FFFFF873FFFFBFBA003FFF840F8786FF;
defparam sp_inst_10.INIT_RAM_2C = 256'hFF000000000000000003004032000003FFFFF831FFFFF9FFF83E006875E040FF;
defparam sp_inst_10.INIT_RAM_2D = 256'hFC00000000000000000216A8F8000007FFE88021FFFF288FF00003E1CBDFC0FF;
defparam sp_inst_10.INIT_RAM_2E = 256'hF000000000000000000A00838E000007FFE20023FFFC0C0603E00946077F003F;
defparam sp_inst_10.INIT_RAM_2F = 256'hC00000000000000004001F000001C003DF000003FFFE08000000B9FFFFFFC20F;
defparam sp_inst_10.INIT_RAM_30 = 256'h00000000000000000067284B9A4180020C008007DFDA1EFEFF85FFF01F007F03;
defparam sp_inst_10.INIT_RAM_31 = 256'h0000000000000000019002C8840180010003C00FF3C13F80E7E7803441F78F00;
defparam sp_inst_10.INIT_RAM_32 = 256'h000000000000000000203A10F80880000003E010C7838001FFE73FF80007C700;
defparam sp_inst_10.INIT_RAM_33 = 256'h0000000000000000000035160803800001F3F0710387C003BF38E0007FFF4000;
defparam sp_inst_10.INIT_RAM_34 = 256'h00000000000000000000C2C1000380000FFDC0E001DDF86BF87FC0007FF98700;
defparam sp_inst_10.INIT_RAM_35 = 256'h00000000000000000020E00E020F80001FFF818002707F3C0FFE0000FFFFFF00;
defparam sp_inst_10.INIT_RAM_36 = 256'h000000000000000000570033DA0F80000FFF02C0001BE3E7FF000001FFF80300;
defparam sp_inst_10.INIT_RAM_37 = 256'h000000000000000000006861932FE00003FF06001BE5CE1EFE18007FFDFA0200;
defparam sp_inst_10.INIT_RAM_38 = 256'h000000000004000000508211C03A500000E30C00101B9FEFC7BC7FE03FC00100;
defparam sp_inst_10.INIT_RAM_39 = 256'h00000000001000000000082E84276A0000608C000E670F41FFFB007F40046000;
defparam sp_inst_10.INIT_RAM_3A = 256'h000000000060000000004007200399400000C80801F0FC078E00007FFFF00800;
defparam sp_inst_10.INIT_RAM_3B = 256'h00000000008000000000011FC0E6C77800000806038770062CE00FFFDCF80000;
defparam sp_inst_10.INIT_RAM_3C = 256'h0000000002000000610000A44217BFFFF000080003EF0E7FFF780FEFFC000000;
defparam sp_inst_10.INIT_RAM_3D = 256'h01000000080000000E00001020C7EFCFF8000800147C2F9FFF8003FE00000000;
defparam sp_inst_10.INIT_RAM_3E = 256'h070000001000100000800000618F5FF3FC0008000001E01FC00C37FFFC200080;
defparam sp_inst_10.INIT_RAM_3F = 256'h1F0000004000000001C081C0405FDBD6DE0000000007C1FFFA00E0FE001800E0;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[30:0],sp_inst_11_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[15],ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b00;
defparam sp_inst_11.BIT_WIDTH = 1;
defparam sp_inst_11.BLK_SEL = 3'b010;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'hFF00000000000000000000000000000000003C003000000700000000000000FF;
defparam sp_inst_11.INIT_RAM_01 = 256'hFF00000000000000000000000000000000001C0020000406C0000000000000FF;
defparam sp_inst_11.INIT_RAM_02 = 256'hFF00000000000000000000000000000000007C004000000F80000000000000FF;
defparam sp_inst_11.INIT_RAM_03 = 256'hFF0000000000000000000000000000000001FE00F800140F00000000000000FF;
defparam sp_inst_11.INIT_RAM_04 = 256'hFF0000000000000000000000000000000000FE00F8001C1E00000000000000FF;
defparam sp_inst_11.INIT_RAM_05 = 256'hFF0000000000000000000000000000000003FE007C003C1C00000000000000FF;
defparam sp_inst_11.INIT_RAM_06 = 256'hFF0000000000000000000000000000000001FE007E00783000000000000000FF;
defparam sp_inst_11.INIT_RAM_07 = 256'hFF0000000000000000000000000000000001FC001F80F06000000000000000FF;
defparam sp_inst_11.INIT_RAM_08 = 256'hFF0000000000000000000000000000000001FE001FFFE04000000000000000FF;
defparam sp_inst_11.INIT_RAM_09 = 256'hFF0000000000000000000000000000000000FC000FFF808000000000000000FF;
defparam sp_inst_11.INIT_RAM_0A = 256'hFF0000000000000000000000000000000001FE0003FF000000000000000000FF;
defparam sp_inst_11.INIT_RAM_0B = 256'hFC0000000000000000000000000000000001FE0000F8000000000000000000FF;
defparam sp_inst_11.INIT_RAM_0C = 256'hF000000000000000000000000000000000007E0000000000000000000000003F;
defparam sp_inst_11.INIT_RAM_0D = 256'hC00000000000000000000000000000000000600000000000000000000000000F;
defparam sp_inst_11.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000003;
defparam sp_inst_11.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_10 = 256'h0000000000000000000000100000000000000000100000000000000000000000;
defparam sp_inst_11.INIT_RAM_11 = 256'h00000000000000000000000000000000000000001A0000000000000000000000;
defparam sp_inst_11.INIT_RAM_12 = 256'h00000000000000000000000000000000000000003FE000000000000000000000;
defparam sp_inst_11.INIT_RAM_13 = 256'h00000000000000000000000000000000000000001FC000000000000000000000;
defparam sp_inst_11.INIT_RAM_14 = 256'h00000000000000000000000000000000000000000F0000000000000000000000;
defparam sp_inst_11.INIT_RAM_15 = 256'h00000000000000000000000000000000000000000D0000000000000000000000;
defparam sp_inst_11.INIT_RAM_16 = 256'h0000000000000000000020000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_17 = 256'h0000000000000000000020000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1B = 256'h0100000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_11.INIT_RAM_1C = 256'h0700000000000000C00000000000000000000000000000000000000000000080;
defparam sp_inst_11.INIT_RAM_1D = 256'h1F000000000000000200000000000000000000000000000000000000000000E0;
defparam sp_inst_11.INIT_RAM_1E = 256'h7F000000000000000200000000000000000000000000000000000000000000F8;
defparam sp_inst_11.INIT_RAM_1F = 256'hFF000000000000000300000000000000000000000000000000000000000000FE;
defparam sp_inst_11.INIT_RAM_20 = 256'hFF000000000000000080000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_21 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_22 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_23 = 256'hFF000000000000000270000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_24 = 256'hFF000000000000000018000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_25 = 256'hFF00000000000000000000000C000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_26 = 256'hFF000000000000000000200178000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_27 = 256'hFF0000000000000000000000F8000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_28 = 256'hFF000000000000000000000000000000000000000000000000000000000000FF;
defparam sp_inst_11.INIT_RAM_29 = 256'hFF00000000000000000000000000000000000000000000000000000000000CFF;
defparam sp_inst_11.INIT_RAM_2A = 256'hFF0000000000000000000000000000000000000000000000000000000007C0FF;
defparam sp_inst_11.INIT_RAM_2B = 256'hFF000000000000000000000000000000000000000000000000000000007801FF;
defparam sp_inst_11.INIT_RAM_2C = 256'hFF0000000000000000000000000000000000000000000000000000000E1F80FF;
defparam sp_inst_11.INIT_RAM_2D = 256'hFC000000000000000000000000000000000000000000000000000000002000FF;
defparam sp_inst_11.INIT_RAM_2E = 256'hF00000000000000000000000000000000000000000000000000000F80080003F;
defparam sp_inst_11.INIT_RAM_2F = 256'hC0000000000000000000000000000000000000000000000000007E000000000F;
defparam sp_inst_11.INIT_RAM_30 = 256'h000000000000000000000000000000000000000020000001007E000000FF8003;
defparam sp_inst_11.INIT_RAM_31 = 256'h00000000000000000000000000000000000000000C00007F00000003FE000000;
defparam sp_inst_11.INIT_RAM_32 = 256'h000000000000000000000000000000000000000F38007FFE0000FFFFFFF80000;
defparam sp_inst_11.INIT_RAM_33 = 256'h000000000000000000000000000000000000000EFC003FFC40FF00000000BF00;
defparam sp_inst_11.INIT_RAM_34 = 256'h000000000000000000000000000000000000001FFE0207940780000000000000;
defparam sp_inst_11.INIT_RAM_35 = 256'h000000000000000000000000000000000000007FFD8F8003F000000000000000;
defparam sp_inst_11.INIT_RAM_36 = 256'h000000000000000000000000000000000000013FFFE400180000000000000000;
defparam sp_inst_11.INIT_RAM_37 = 256'h00000000000000000000000000000000000001FFE41A000101E0000000000000;
defparam sp_inst_11.INIT_RAM_38 = 256'h00000000000000000000000000000000000003FFEFE000103803FFFFC0000000;
defparam sp_inst_11.INIT_RAM_39 = 256'h00000000000000000000000000000000000003FFF18000BE00040000BFFF8000;
defparam sp_inst_11.INIT_RAM_3A = 256'h00000000000000000000000000000000000007F7FE0003F87000000000000700;
defparam sp_inst_11.INIT_RAM_3B = 256'h00000000000000000000000000000000000007F9FC000FF9FF00000000000000;
defparam sp_inst_11.INIT_RAM_3C = 256'h00000000000000000000000000000000000007FFFC00F1800007FFF000000000;
defparam sp_inst_11.INIT_RAM_3D = 256'h01000000000000000000000000000030000007FFEB83D00000000001F8000000;
defparam sp_inst_11.INIT_RAM_3E = 256'h0700000000000000000000000000000C000007FFFFFE00003FF0000003C00080;
defparam sp_inst_11.INIT_RAM_3F = 256'h1F00000000000000000000000000002920000FFFFFF8000000001F00000700E0;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[29:0],sp_inst_12_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[15],ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b00;
defparam sp_inst_12.BIT_WIDTH = 2;
defparam sp_inst_12.BLK_SEL = 3'b110;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'hCF3C4450422FFA828C55E4D4F56A5BEABFE903EBFF56238BD2E9AA599135FFC0;
defparam sp_inst_12.INIT_RAM_01 = 256'h3FFF555555555557D55556AA556AA5550085ED58906FE3F3EDACEC0A36F5BD13;
defparam sp_inst_12.INIT_RAM_02 = 256'h30430040021AA6940D4FBE043C0C53EA540E8C030EC309ACEB69D95A95D0FFFC;
defparam sp_inst_12.INIT_RAM_03 = 256'hFFFF55555555555955556EBA959655550041E15E5555CAF3AA8FE4C70848F231;
defparam sp_inst_12.INIT_RAM_04 = 256'hC01880000BDAAA911400316BEFEAACF98AACA56AABFC3CFFC043FD7A6BACFFFF;
defparam sp_inst_12.INIT_RAM_05 = 256'hFFFF5555555555355555596A95551555054554594659AFB2ABAB3FA5B213B207;
defparam sp_inst_12.INIT_RAM_06 = 256'h00D53910540659A56B00505BCFA951A8B0329FBAAA68143D8C143BAC3A03FFFF;
defparam sp_inst_12.INIT_RAM_07 = 256'hFFFF555555555555555955AA95544450001555655556BF8EAA611B943B56B41C;
defparam sp_inst_12.INIT_RAM_08 = 256'h0F55411977800914E36AC1AAFFA501AA4157B45BBEAEACD000100EBA6C0DFFFF;
defparam sp_inst_12.INIT_RAM_09 = 256'hFFFF555555554155555555599500441400555955559A6FFA4D615B559059D8D3;
defparam sp_inst_12.INIT_RAM_0A = 256'hC1559650CCD7B0CFCDE9AC0F5335268A40EA6658BE95570B33C4FE5BFCC1FFFF;
defparam sp_inst_12.INIT_RAM_0B = 256'hFFFF55555554955555555556A9505404056565555A5AA56AA9A919FAA027ACCF;
defparam sp_inst_12.INIT_RAM_0C = 256'hCD55633951309BDAB3FC3F0833F15AA29F95AA3CD4F56EAFC3C0EA6ABC00FFFF;
defparam sp_inst_12.INIT_RAM_0D = 256'hFFFF5555555D55555555559AA9510104155999955556A9AAD922A043829FFFEF;
defparam sp_inst_12.INIT_RAM_0E = 256'hE00555D352AFEB0AAFE9AA57AF915BA500856BC02A1BFAFB9104A5E56BFFFFFF;
defparam sp_inst_12.INIT_RAM_0F = 256'hFFFF55555565555555599556AA510565969AA6AAAA9A96BA98BFF0511172ABBF;
defparam sp_inst_12.INIT_RAM_10 = 256'h8CC456585567FFFD6850D468001355AA3BBAEC501728097ABB0655B26F0CFFFF;
defparam sp_inst_12.INIT_RAM_11 = 256'hFFFF55555055555555955556695111556659AAAAAA6957AA6AB54298103893FA;
defparam sp_inst_12.INIT_RAM_12 = 256'h3C00E41E5025AFEA9AAFF559030609938D9BFF8CC896C9CC12F950783DF9FFFF;
defparam sp_inst_12.INIT_RAM_13 = 256'hFFFF55555955555555555555AEE54154555A9AAAAA9556A580264E510F546B7B;
defparam sp_inst_12.INIT_RAM_14 = 256'hF30D7C090055AAAB6A6AA996B006FFBEBC03154E9F9425C3455D956FAB01FFFF;
defparam sp_inst_12.INIT_RAM_15 = 256'hFFFF5555A555555555556A66FE95551166969AAA5699591AC65A57D7D91099AF;
defparam sp_inst_12.INIT_RAM_16 = 256'hCF3A78A5C01565AFF5AAEF5140556AB4AB190512AABEA5ABB4E955AC0190FFFF;
defparam sp_inst_12.INIT_RAM_17 = 256'hFFFF5554555555555555565EBBA55546969AAAA9BAA651AF15554FEA9BDF5A7F;
defparam sp_inst_12.INIT_RAM_18 = 256'hEFEEEB84FF74357A7AA9A9555159A64093C214027C676F315715555B3111FFFF;
defparam sp_inst_12.INIT_RAM_19 = 256'hFFFF555055555555555555555BFA9A66A9AAAABBFEE56AAB54733F66BE40AABF;
defparam sp_inst_12.INIT_RAM_1A = 256'h6EAAF682AAFC29566896950001A943CFEE84401E5DD7D381099659AAF409FFFF;
defparam sp_inst_12.INIT_RAM_1B = 256'hFFFF551555555555555555555BFA95996AAAAAFAAA55AAA80CCECE562016A4AE;
defparam sp_inst_12.INIT_RAM_1C = 256'h2A3AE502AAAB345118145004415A44F02CB9901925572ECA6A5596BFB008FFFF;
defparam sp_inst_12.INIT_RAM_1D = 256'hFFFF555555555555555555555AFEA6AA9AAA6FEA5551AAAF134AC03A9C56A166;
defparam sp_inst_12.INIT_RAM_1E = 256'hA669950E5A6AA4F0F783000156A59CF31015554272A800109969D95FEF03FFFF;
defparam sp_inst_12.INIT_RAM_1F = 256'hFFF07D55555555555555554556AEAA5AAFEAFEA9655A6AB7330ED54171764748;
defparam sp_inst_12.INIT_RAM_20 = 256'h59A9140A999AB7ECFFCFC0555559553AC5FA54C00F112AFCADAA68A6AAFA0FFF;
defparam sp_inst_12.INIT_RAM_21 = 256'hFF00D555555555555555555555BBA65AAAAFF9A999AAAE260C1C555584C04015;
defparam sp_inst_12.INIT_RAM_22 = 256'h3AA9573956597BAFFC031556A95026F98111AA530670EBBBEBFA5BC76B3E00FF;
defparam sp_inst_12.INIT_RAM_23 = 256'hF0005555555555555555555555AEA95AAA6EA5B9A5693639F55995550CCF5556;
defparam sp_inst_12.INIT_RAM_24 = 256'hA56917395A6ABAECC01555559654FAABFD45479505C83FFE8FE591668B1F000F;
defparam sp_inst_12.INIT_RAM_25 = 256'h000055555555555555555555555ABAA5A6959B9EAAAB5BCBD56A534BB3415545;
defparam sp_inst_12.INIT_RAM_26 = 256'hA85513FAAA6FE3EF00555A955553F9980C5C65101555149BB2F56EEEB4C30000;
defparam sp_inst_12.INIT_RAM_27 = 256'h000055555555555555555555556EFAAA9959BD3AAA2588EA5400F6AE80525895;
defparam sp_inst_12.INIT_RAM_28 = 256'h9455FEBA9EACEF00C55AAAA9150FFFBF545FB996424D44E9F80259AEB34F0000;
defparam sp_inst_12.INIT_RAM_29 = 256'h000055555555555555555555557AEBEEA595DEA5A254FD56100AE5AAC4446356;
defparam sp_inst_12.INIT_RAM_2A = 256'h9450FA8FABFCE3F0D56AAAA9503E7F00F156A83C41515F556B4FEABFBFF10000;
defparam sp_inst_12.INIT_RAM_2B = 256'h000055555555555555555555565BAABAA559A544112DD944980F3CF315315046;
defparam sp_inst_12.INIT_RAM_2C = 256'h540CEA8FA733C33C019AAAAA5432FC10FB012AF7F8001495FFD0BB9BCDAF0000;
defparam sp_inst_12.INIT_RAM_2D = 256'h000055555555555555555555556F96BBA9A6558D546C5A1595F0C00010EC4355;
defparam sp_inst_12.INIT_RAM_2E = 256'h400F3B8FA0CCC17716BAAA6953F8F1065705CE92C30E1356EB42A58FAC130000;
defparam sp_inst_12.INIT_RAM_2F = 256'h00005555555555555555555555AA966BAAE9585557D542114D7C002301AC5C15;
defparam sp_inst_12.INIT_RAM_30 = 256'h3F0C3B83F00F011511FF955543ABD1A6B10030BAAB0C9565BBF0F556ACFF0000;
defparam sp_inst_12.INIT_RAM_31 = 256'h000055555555555555555555569AA6AAE2AB36A50A65514345AECB83F3E03C10;
defparam sp_inst_12.INIT_RAM_32 = 256'hF00C23C300104686516B95400EBBB35554003F4BBFCF94185B01FE556FBE0000;
defparam sp_inst_12.INIT_RAM_33 = 256'h0000555555555555555555595966AAAAFE929AA5B958055D1507286FF3FDF004;
defparam sp_inst_12.INIT_RAM_34 = 256'hC0000000C0554595545A9400FBFFEE1595525F1430CEA45693303F3AB33B0000;
defparam sp_inst_12.INIT_RAM_35 = 256'h0000559555955555555555559555BAACA4EAAB4EA9D2A4F5559A507CC3000003;
defparam sp_inst_12.INIT_RAM_36 = 256'h00055C51D11596A99455500FEAB0FA4DA550F4E753FB596B17FF3EB9EB3B0000;
defparam sp_inst_12.INIT_RAM_37 = 256'h0000555555655555555555555556A9DBD6AAAB2BEE069B5554357EA27F00C003;
defparam sp_inst_12.INIT_RAM_38 = 256'h001440D1165655AD510150EEABFF12966950CDCA572955959FC3AD5AE6BE0000;
defparam sp_inst_12.INIT_RAM_39 = 256'h00005595555A55955555556565A9A547EEAAA3BAD8EA415669C5F5A83F0F0000;
defparam sp_inst_12.INIT_RAM_3A = 256'h41554C112A6565BD544503AAAAC044F8D625AB412AA455ABCAAABAAAEAAA0000;
defparam sp_inst_12.INIT_RAM_3B = 256'h000055555555E555555555556AAAB08FFBADFA99D6BB5695B742E944BF2F0000;
defparam sp_inst_12.INIT_RAM_3C = 256'h55554CC166559459555030AABEED6A394A266D5FE55A554F38EAE97A96AA0000;
defparam sp_inst_12.INIT_RAM_3D = 256'h0000556555555B55555555559BA42ABEE3B2AE43DFE7AAA9840EE5BABBEFC000;
defparam sp_inst_12.INIT_RAM_3E = 256'h155510D19555555A5513FB2AECFB3FA2878B25CD541666DFBF66BEDC69AA0000;
defparam sp_inst_12.INIT_RAM_3F = 256'h000355555555557355555556CB5EEAAA0F12D6F8FF9EAAA711A8552EAEAEF001;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[29:0],sp_inst_13_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({ad[15],ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b00;
defparam sp_inst_13.BIT_WIDTH = 2;
defparam sp_inst_13.BLK_SEL = 3'b110;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'h6595000001AAAAAAA6AA5515000555555555540000554415540000001A80FFC0;
defparam sp_inst_13.INIT_RAM_01 = 256'h3FFF0000000000000000000000000000000000010000040400010150450556A9;
defparam sp_inst_13.INIT_RAM_02 = 256'h9AA9400001AAAAAAA6A555554156A955555011545014500100550000001AFFFC;
defparam sp_inst_13.INIT_RAM_03 = 256'hFFFF00000000000400000000000000000000000000001004001004105155599A;
defparam sp_inst_13.INIT_RAM_04 = 256'h6AAA5000016AAAAAAAAA9555555556AA5001000000014100155401400001FFFF;
defparam sp_inst_13.INIT_RAM_05 = 256'hFFFF0000000000400000000000000000000000000000000400000000045559A9;
defparam sp_inst_13.INIT_RAM_06 = 256'hAA6A900001AAAAAA95AAA95565555556AFE9500000015541515540014054FFFF;
defparam sp_inst_13.INIT_RAM_07 = 256'hFFFF0000000001000000000000000000000000000000001000000000005556A6;
defparam sp_inst_13.INIT_RAM_08 = 256'hA5AAA500056AAAAA59556A55555555555555A90000000115555550000151FFFF;
defparam sp_inst_13.INIT_RAM_09 = 256'hFFFF000000001400000000000000000000000000000000001000000005555659;
defparam sp_inst_13.INIT_RAM_0A = 256'h6AAAA90412695A65655556A554455AA55500006A00000050441500000115FFFF;
defparam sp_inst_13.INIT_RAM_0B = 256'hFFFF000000004000000000000000000000000000000000000000000005555665;
defparam sp_inst_13.INIT_RAM_0C = 256'h66AAA940559A5555595695A54405555AA400004169000000141500000155FFFF;
defparam sp_inst_13.INIT_RAM_0D = 256'hFFFF000000010000000000000000000000000000000000000004055415555555;
defparam sp_inst_13.INIT_RAM_0E = 256'h5AAAAA54555555A55555555401555555556A401541A40000555500000000FFFF;
defparam sp_inst_13.INIT_RAM_0F = 256'hFFFF000000100000000000000000000000000000000000000000055555595555;
defparam sp_inst_13.INIT_RAM_10 = 256'h666AAA955555555556AA555555595555400016955441A540005000040051FFFF;
defparam sp_inst_13.INIT_RAM_11 = 256'hFFFF000001000000000000000000000000000000000000000005555555555955;
defparam sp_inst_13.INIT_RAM_12 = 256'h96AA5A9555555555555555555455A5541000001655001651540000014100FFFF;
defparam sp_inst_13.INIT_RAM_13 = 256'hFFFF000004000000000000000000000000000000000000001555555550555555;
defparam sp_inst_13.INIT_RAM_14 = 256'h59A556A55555555555555555455555400154555015554019555000000055FFFF;
defparam sp_inst_13.INIT_RAM_15 = 256'hFFFF000000000000000000000000000000000000000000001555541400555555;
defparam sp_inst_13.INIT_RAM_16 = 256'h659556551555555555555555555555550055555400500000550000015555FFFF;
defparam sp_inst_13.INIT_RAM_17 = 256'hFFFF000100000000000000000000000000000000000000005555500000105555;
defparam sp_inst_13.INIT_RAM_18 = 256'h555555150045455555555555555555555415555541554045554000004555FFFF;
defparam sp_inst_13.INIT_RAM_19 = 256'hFFFF000400000000000000000000000000000000000000005544400000555555;
defparam sp_inst_13.INIT_RAM_1A = 256'h555555140001455555555555555554100155555055001415501400000555FFFF;
defparam sp_inst_13.INIT_RAM_1B = 256'hFFFF004000000000000000000000000000000000000000015110100045555555;
defparam sp_inst_13.INIT_RAM_1C = 256'h555555540000455555555555555555054155555555544115400140000555FFFF;
defparam sp_inst_13.INIT_RAM_1D = 256'hFFFF010000000000000000000000000000000000000000004450154051555555;
defparam sp_inst_13.INIT_RAM_1E = 256'h555555500000010504145555555551045555555545555555500014000054FFFF;
defparam sp_inst_13.INIT_RAM_1F = 256'hFFF0000000000000000000000000000000000000000000040450155545455455;
defparam sp_inst_13.INIT_RAM_20 = 256'h5555555000000001001015555555554015055515505540010000014000000FFF;
defparam sp_inst_13.INIT_RAM_21 = 256'hFF00000000000000000000000000000000000000000001405151555555155555;
defparam sp_inst_13.INIT_RAM_22 = 256'h55555440000000000154555555554000155555545405000000000014004000FF;
defparam sp_inst_13.INIT_RAM_23 = 256'hF000000000000000000000000000000000000000000054410555555551105555;
defparam sp_inst_13.INIT_RAM_24 = 256'h555554400000000115555555555500000155545555114000100000005050000F;
defparam sp_inst_13.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000505101555545004555555;
defparam sp_inst_13.INIT_RAM_26 = 256'h5555540000000400555555555554000151515555555555000400000005140000;
defparam sp_inst_13.INIT_RAM_27 = 256'h0000000000000000000000000000000000000040009021005555000015555515;
defparam sp_inst_13.INIT_RAM_28 = 256'h5555000000010055155555555550000055500555555155000154000004500000;
defparam sp_inst_13.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000180200055550040015555455;
defparam sp_inst_13.INIT_RAM_2A = 256'h5555001000010405155555555540005505540141555550000050000000050000;
defparam sp_inst_13.INIT_RAM_2B = 256'h0000000000000000000000000000000000000002401400250150510455455555;
defparam sp_inst_13.INIT_RAM_2C = 256'h5551001000441441555555555544015500554000015555000015000011000000;
defparam sp_inst_13.INIT_RAM_2D = 256'h0000000000000000000000000000000000000020008000900505555555015455;
defparam sp_inst_13.INIT_RAM_2E = 256'h5550401005111544555555555401055554551004145054000054001001540000;
defparam sp_inst_13.INIT_RAM_2F = 256'h0000000000000000000000000000000000000600080005002002555455015155;
defparam sp_inst_13.INIT_RAM_30 = 256'h4051401405505555555555555400155545554500005100000005000001000000;
defparam sp_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000004008000900020014004105404054155;
defparam sp_inst_13.INIT_RAM_32 = 256'h0551441455555555555555555000045555554050001000000055000000000000;
defparam sp_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000180002000280040020415004010555;
defparam sp_inst_13.INIT_RAM_34 = 256'h1555555515555555555555550000005555545055451000000045404004400000;
defparam sp_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000106000020001800400044054114555554;
defparam sp_inst_13.INIT_RAM_36 = 256'h5555515515555555555555500005005155550514540000005400400000400000;
defparam sp_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000001050000080016001000210110440551554;
defparam sp_inst_13.INIT_RAM_38 = 256'h5555551555555555555555000000541455551115544000000014000000000000;
defparam sp_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000016400000800120024000440440140505555;
defparam sp_inst_13.INIT_RAM_3A = 256'h5555515555555555555554000015550515555455400000001000000000000000;
defparam sp_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000191000001005180080000401001500405555;
defparam sp_inst_13.INIT_RAM_3C = 256'h5555511555555555555545000001554555455550000000104100000000000000;
defparam sp_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000006400004004054500500006000000000001555;
defparam sp_inst_13.INIT_RAM_3E = 256'h5555551555555555555400400100555555505510000000000000000100000000;
defparam sp_inst_13.INIT_RAM_3F = 256'h0003000000000004000000001550000050481406002000018041004000000555;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[27:0],sp_inst_14_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[11:0],gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:0]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b00;
defparam sp_inst_14.BIT_WIDTH = 4;
defparam sp_inst_14.BLK_SEL = 3'b001;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h55356654444243110110110122333433222322313222224422221122F0000000;
defparam sp_inst_14.INIT_RAM_01 = 256'h4555554545444555656554554555555555543442222122433423444445666665;
defparam sp_inst_14.INIT_RAM_02 = 256'h2324484432344934443652222223327321261322211232121222222233333344;
defparam sp_inst_14.INIT_RAM_03 = 256'h00000FFF11111111111111111111111112445444445677221224321122212233;
defparam sp_inst_14.INIT_RAM_04 = 256'h55436665533213200011111123243344555332331232322333223121FFF00000;
defparam sp_inst_14.INIT_RAM_05 = 256'h4555555554545455655544554554555555543342122222233433343563567656;
defparam sp_inst_14.INIT_RAM_06 = 256'h2145734433374343226512222322282215423411121512111222212322233344;
defparam sp_inst_14.INIT_RAM_07 = 256'h000FFFFF11111111111111111111111111110101124301112342221222221312;
defparam sp_inst_14.INIT_RAM_08 = 256'h44444556545110110010010232243433332434221223322212322221FFFFF000;
defparam sp_inst_14.INIT_RAM_09 = 256'h3454455544555444555544444444454555442331213223334435423357454654;
defparam sp_inst_14.INIT_RAM_0A = 256'h5345333335733333482323333222912262232223223121212211112221322333;
defparam sp_inst_14.INIT_RAM_0B = 256'h0FFFFFFF11111111111111111111111111111111101112343232222222212223;
defparam sp_inst_14.INIT_RAM_0C = 256'h44353433423210010111123323333244444222321211133343222221FFFFFFF0;
defparam sp_inst_14.INIT_RAM_0D = 256'h3344445445454545555545444444454455442222222222445564452435754545;
defparam sp_inst_14.INIT_RAM_0E = 256'h2452333284433334733344421228123522262332223321112111111112222333;
defparam sp_inst_14.INIT_RAM_0F = 256'hFFFFFFFF11111111111111111111111111111111111124333321122211124531;
defparam sp_inst_14.INIT_RAM_10 = 256'h44433132011212112112123224423433324311122112232311222221FFFFFFFF;
defparam sp_inst_14.INIT_RAM_11 = 256'h3333454444444455555444444444444454333222122223234776555423364442;
defparam sp_inst_14.INIT_RAM_12 = 256'h5212225632424366333434322383243332733233243221221111111122222233;
defparam sp_inst_14.INIT_RAM_13 = 256'hFFFFFFFF11111111111111111111110111111111112322322322222443211121;
defparam sp_inst_14.INIT_RAM_14 = 256'h23232211010111111112323433332343123233223432333222222221FFFFFFFF;
defparam sp_inst_14.INIT_RAM_15 = 256'h1333333444444454545444444443344444312323122221423566755431325432;
defparam sp_inst_14.INIT_RAM_16 = 256'h2111181222343734333452323744532227322322432222211111111111221122;
defparam sp_inst_14.INIT_RAM_17 = 256'hFFFFFFFF11111111111111111111110110111111311112223454221112211215;
defparam sp_inst_14.INIT_RAM_18 = 256'h21222111111111111122223343322133201244221433333331111111FFFFFFFF;
defparam sp_inst_14.INIT_RAM_19 = 256'h1223323343334444544444444443334433211243212222221355665463243342;
defparam sp_inst_14.INIT_RAM_1A = 256'h1213513222237322343443347445333364233322332321212111121111111121;
defparam sp_inst_14.INIT_RAM_1B = 256'hFFFFFFFF11111111111111111111111101111121111134432222221111112161;
defparam sp_inst_14.INIT_RAM_1C = 256'h10101112111101111123243343431222331112332123233322311211FFFFFFFF;
defparam sp_inst_14.INIT_RAM_1D = 256'h1122211432233243444433334343323321212113313224322135364654022213;
defparam sp_inst_14.INIT_RAM_1E = 256'h1182222222362333443344374554333433332333213232232211211112111111;
defparam sp_inst_14.INIT_RAM_1F = 256'hFFFFFFFF11111211111111111111111111111002432222222222211111121612;
defparam sp_inst_14.INIT_RAM_20 = 256'h10110021211111211113444222232233211112232122333332222311FFFFFFFF;
defparam sp_inst_14.INIT_RAM_21 = 256'h1121114322222333333433334333223322222123322244433322344554311123;
defparam sp_inst_14.INIT_RAM_22 = 256'h6212121214643234433344835333333533434343333323323222221121211111;
defparam sp_inst_14.INIT_RAM_23 = 256'hFFFFFFFF21111111111111111111111111113211111222122222211112225322;
defparam sp_inst_14.INIT_RAM_24 = 256'h11111111111111112422454422242222321322322322122242213201FFFFFFFF;
defparam sp_inst_14.INIT_RAM_25 = 256'h1211122222222232333322333322212322222313352334533423333463501112;
defparam sp_inst_14.INIT_RAM_26 = 256'h1211112145323333323337253333325334443343333232322122221112122111;
defparam sp_inst_14.INIT_RAM_27 = 256'hFFFFFFFF21211111111111111111111112110111111112222222211222243217;
defparam sp_inst_14.INIT_RAM_28 = 256'h11111121111112343442333342325313323212122233433323311122FFFFFFFF;
defparam sp_inst_14.INIT_RAM_29 = 256'h1211222222222222222232233222222123424322343244433323343343311110;
defparam sp_inst_14.INIT_RAM_2A = 256'h1111111632243333233374543334313443234433332323331222112322121111;
defparam sp_inst_14.INIT_RAM_2B = 256'hFFFFFFFF11121111111111111011110111111111111112222222222226232341;
defparam sp_inst_14.INIT_RAM_2C = 256'h21111113121112253243223334433300211231212324433323332111FFFFFFFF;
defparam sp_inst_14.INIT_RAM_2D = 256'h1222232221222222222233222222431122434422244234423222322334111021;
defparam sp_inst_14.INIT_RAM_2E = 256'h1111116321443332222544213321253213434334331333312222123121222111;
defparam sp_inst_14.INIT_RAM_2F = 256'hFFFFFFFF11111111111111111111111111110101100112222222222262334412;
defparam sp_inst_14.INIT_RAM_30 = 256'h21112212211111233314322433422233112121121243243312332311FFFFFFFF;
defparam sp_inst_14.INIT_RAM_31 = 256'h1222222222222323233233223222231112143422222222113211212123121111;
defparam sp_inst_14.INIT_RAM_32 = 256'h1212171113233322214622210111111323233433333322123221232221222222;
defparam sp_inst_14.INIT_RAM_33 = 256'hFFFFFFFF11121111111111111110111101001111111133222333326433353111;
defparam sp_inst_14.INIT_RAM_34 = 256'h21111222231221122311422254453212321123223323333443201341FFFFFFFF;
defparam sp_inst_14.INIT_RAM_35 = 256'h2232222322222323233233223222132001132431110211101121201121311211;
defparam sp_inst_14.INIT_RAM_36 = 256'h1111511111222222155021011112522222333333332222222222323222122222;
defparam sp_inst_14.INIT_RAM_37 = 256'hFFFFFFFF11111211111111111100011001011111112233232333553433422322;
defparam sp_inst_14.INIT_RAM_38 = 256'h11111222222111324331232433434243322111222344334344211112FFFFFFFF;
defparam sp_inst_14.INIT_RAM_39 = 256'h3233322333222333233233323322132010122331011111000002200221211111;
defparam sp_inst_14.INIT_RAM_3A = 256'h1115111122112222252111111221111111323322221222232223233232223233;
defparam sp_inst_14.INIT_RAM_3B = 256'hFFFFFFFF11111111111111111101000001101111123333332336233333423221;
defparam sp_inst_14.INIT_RAM_3C = 256'h11012222222343133524221132231323312212222223443312211111FFFFFFFF;
defparam sp_inst_14.INIT_RAM_3D = 256'h3333322323312323233233332312122000012221111111111101311122111122;
defparam sp_inst_14.INIT_RAM_3E = 256'h1341111221112112632121112114111112211211122311223222343322232233;
defparam sp_inst_14.INIT_RAM_3F = 256'hFFFFFFFF11111111111111111101111110010001122222223513334434443311;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce_w)
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(sp_inst_12_dout[0]),
  .I1(sp_inst_14_dout[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(sp_inst_0_dout[0]),
  .I1(sp_inst_1_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(sp_inst_8_dout[0]),
  .I1(mux_o_8),
  .S0(dff_q_1)
);
MUX2 mux_inst_11 (
  .O(dout[0]),
  .I0(mux_o_9),
  .I1(mux_o_10),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(sp_inst_12_dout[1]),
  .I1(sp_inst_14_dout[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sp_inst_2_dout[1]),
  .I1(sp_inst_3_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(sp_inst_9_dout[1]),
  .I1(mux_o_20),
  .S0(dff_q_1)
);
MUX2 mux_inst_23 (
  .O(dout[1]),
  .I0(mux_o_21),
  .I1(mux_o_22),
  .S0(dff_q_0)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(sp_inst_13_dout[2]),
  .I1(sp_inst_14_dout[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(sp_inst_4_dout[2]),
  .I1(sp_inst_5_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(sp_inst_10_dout[2]),
  .I1(mux_o_32),
  .S0(dff_q_1)
);
MUX2 mux_inst_35 (
  .O(dout[2]),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sp_inst_13_dout[3]),
  .I1(sp_inst_14_dout[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(sp_inst_6_dout[3]),
  .I1(sp_inst_7_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(sp_inst_11_dout[3]),
  .I1(mux_o_44),
  .S0(dff_q_1)
);
MUX2 mux_inst_47 (
  .O(dout[3]),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(dff_q_0)
);
endmodule //Gowin_SP
