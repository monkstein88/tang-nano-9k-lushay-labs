// In this article we will be taking a look at generating pseudo-random numbers using an LFSR (Linear Feedback Shift Register) and look at how one can be used as part of a larger application.
//
// The LFSR
// An LFSR is a shift register like we have seen in previous articles, except that the bits besides shifting are also affected by the other bits in the register - this effect is what is referred 
// to as the feedback.
//
// There are multiple variations of LFSR but in this article we will be focusing on the most basic type the Fibonacci LFSR. In this type of LFSR the feedback only affects the first bit. So all 
// bits get shifted up and the least significant bit is generated using the feedback of the current registers bits.
// 
// A basic example of a 5-bit LFSR:
//
//                                /-----|| 
//                               /      ||<----------------------+
//               +--------------{  XOR  ||                       |
//               |               \      ||<--+                   |
//               |                \-----||   |                   |
//               |                           |                   |
//               |                           |                   |
//               |                 +-----+---*--+------+-----+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |  B3 |  B4  |-------| >
//                 LSFR INPUT BIT  |     |      |      |     |      |       |/
//                                 +-----+------+------+-----+------+
//                                   LSb                        MSb
//                                     
// So in the example above on each clock cycle B4 is the output bit b0-b3 get shifted up and a new bit is generated by XOR-ing bit 4 and bit 1 this new bit gets inserted into b0.
//
// The bits we choose for our feedback are called "taps", and not every arrangement of taps are good options. Since our new bit is generated by XOR-ing bits, if all bits were zero the system 
// would be stuck in the zero state. XOR can be thought of as returning 1 if the number of 1s being XOR-ed is odd. Since all zeroes has zero 1s and shifting will just keep inputting a new zero
// we never get out of this state.
//
// Another thing to consider, the entire equation is only based on the current state of the register there is no other state being used in the calculation, so as soon as the register rolls 
// back to a number it already was on that will create a cycle. For example if we have an LFSR generating numbers from 1-16 but has an initial cycle of: 1, 4, 7, 14, 3, 5, 7, 14, 3, 5, 7
//
// You can see that as soon as we had two ways of getting to 7 (both 4 generated a 7 as the next number and also a 5) we get stuck in a loop between the two numbers. All further cycles will just
// go between 7, 14, 3, 5 in an endless cycle.
//
// The problem with these short cycles is that the LFSR can no longer generate any number in the range. If I have a 6-sided dice that can only be a 2 or a 4 it wouldn't really be considered a 
// fair dice in the realm of numbers 1-6 as the probabilities for each number are not the same.
//
// So when choosing taps we want to choose something that:
// 1. Never generates all zeroes
// 2. Generates a sequence that goes through all possible numbers
//
// Luckily for us, we do not have to manually calculate optimal taps instead there are pre-calculated tables for max length taps. For example this site here has a precompiled list of max-length 
// taps for LFSRs with 4-64 bits.
//
// For example opening the file for 5-bit LFSRs like in the example above has the following options:
// 0x12
// 0x14
// 0x17
// 0x1B
// 0x1D
// 0x1E
//
// Each of these is an optional tap set. The example above used the 12 option, these numbers are in hex, but converting 12 hex to binary provides:
// 0b10010
//
// Least significant bit to least significant bit, this means take bits index 1 and index 4 for the feedback and leave out index 0,2 and 3 like in this image:
//
//                                /-----|| 
//                               /      ||<----------------------+
//               +--------------{  XOR  ||                       |
//               |               \      ||<--+                   |
//               |                \-----||   |                   |
//               |                           |                   |
//               |                           |                   |
//               |                 +-----+---*--+------+-----+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |  B3 |  B4  |-------| >
//                 LSFR INPUT BIT  |     |      |      |     |      |       |/
//                                 +-----+------+------+-----+------+
//                                   LSb                        MSb
//
// But any of these options would produce a max-length sequence. Now that we have something that can generate a complete sequence of all numbers let us talk a little about the "random" part.
//
//
// Pseudo Random
//
// The LFSR produces a sequence which includes all the possible options, but that doesn't necessarily make it "random". For example if we are talking about a 3-bit LFSR, we can get all the numbers
// 1-7, but a 3-bit counter also produces all the numbers from 1-7 but it would hardly be random.
//
// Taking a look at a counter's sequence:  
// 1,2,3,4,5,6,7
//
// All numbers in this sequence have the same number of occurrences, but each number is just the previous number plus 1 making it to obvious of a relationship for us to call it unpredictable 
// or random.
//
// Now like with a deck of cards, the way can randomize the output is by shuffling. So let's shuffle this group of numbers into the following for example:
// 7, 6, 4, 1, 2, 5, 3
//
// One can now say that the sequence is random, because the order in which the numbers come out are no longer related to previous elements. The sequence is still not perfect as there are no duplicates,
// for example with rolling a dice I can roll a 4 and then roll another 4 before going through all the other options. But we can at least say it is as random as a deck of cards being randomly shuffled.
// 
// The problem with this solution is it requires something else to randomly shuffle the elements for it to really be random and it is hardware intensive to implement. To create such a system we would 
// need to store each number of the sequence kind of like a 1-time pad so for example with a 32-bit LFSR we would need to store 2^32 -1 numbers over 4-billion 32-bit numbers or about 16GB of storage 
// for 1 sequence, and we would even want sequences much longer then this.
//
// So an LFSR is somewhere in-between a real shuffled sequence to a sequence with an obvious relation like a counter. The LFSR - when the taps are chosen correctly - produces all the numbers (except 0)
// in a sequence shuffled based on a non-obvious relation.
//
//
//                                /-----||      
//                               /      ||<---------+
//               +--------------{  XOR  ||          |
//               |               \      ||<--+      |
//               |                \-----||   |      |
//               |                           |      |
//               |                           |      |
//               |                 +-----+---*--+---*--+       |\  LSFR OUTPUT BIT
//               +---------------->|  B0 |  B1  |  B2  |-------| >
//                 LSFR INPUT BIT  |     |      |      |       |/
//                                 +-----+------+------+
//                                   LSb           MSb
//
// Starting with the seed value (initial value) of 1, let's the sequence given by this shift register will be:
// binary  | decimal
//  001    | 1
//  011    | 3
//  111    | 7
//  110    | 6
//  101    | 5
//  010    | 2
//  100    | 4
//  001    | 1
//
// Looking at this sequence you can see that we go through all the numbers before reaching back to 1 and that the sequence is shuffled. The reason we call this "pseudo-random" and not random is because 
// there is a correlation between them, it can be said that the function for the first bit is:
// b0 = b1 xor b2
// and that for the other bits the equation is simply:
// b_i = b_(i-1)
//
// As each bit is simply shifted up. Since there is a correlation between the previous state and the next state with enough of the sequences outputs one could solve some math equations and work out which 
// taps were chosen being able to predict future numbers in the sequence.
//
// So it's not unpredictable, but the order has no meaningful meaning so we can say it is shuffled. With that said there are some things we can do to make it even better.
//
// The first thing is to make the LFSR larger then the number we are using. For example if we need a 4-bit number and we use instead a 5-bit LFSR taking 4 bits at a time, we essentially doubled the number
// of times each number comes up allowing our sequence to have streaks of the same number like we mentioned that dice rolls have. We also get the ability to get 0 as a number, all the bits of an LFSR 
// cannot equal zero but if you are reading only some of the bits then they can all equal zero.
//
// In reality you usually want the LFSR to be much bigger (not just by one bit) and use a relatively small number of bits. Another way to make it better is to not reuse the same bits and to skip bits 
// in-between numbers.
//
// Each shift of the register you only get 1 new "random" bit. All the other bits are just shifted over which is like doubling. So in the case of the 3-bit LFSR if you wait 3-bits before taking another
// number then all of the new numbers 3-bits are completely unrelated to the bits of the previous number making it more random.
//
// Finally if you let the LFSR run in the background essentially skipping generated bits and then let random actions like when a user pressed a button decide when to read the next number you are 
// essentially adding in random like when shuffling bringing it closer to real random.
//
// I think that is enough theory though let's get into building this.
//
//
// Generalizing the LFSR Module
// The difference between all LFSRs of this type (fibonacci / external LFSRs) is the size of the register (num bits) the tap configuration, and some would say the initial seed.
// Changing the seed doesn't change the sequence, it just changes where you start in the sequence, but we can say that this is another difference.
// Other then that we still just need to create a register shift the bits over and calculate the new bit based on the taps chosen.
// Let's create a file called lfsr.v with a module accepting these as parameters:

`default_nettype none 

module lfsr 
#(
  parameter SEED = 5'd1,
  parameter TAPS = 5'h1B,
  parameter NUM_BITS = 5
)
(
  input  wire clk,
  output reg  randomBit 
);
  reg [NUM_BITS-1:0] sr = SEED; //  create a register of the desired size holding our seed value as it's initial value
  wire finalFeedback; // a wire which will hold the feedback after the feedback calculation (XORs). 
  
  always_ff@(posedge clk) begin   // The calculation each clock cycle:
    sr <= {sr[NUM_BITS-2:0], finalFeedback}; // shifting all the bits up 1 and putting our feedback bit into b0.
    randomBit <= sr[NUM_BITS-1]; // output bit
  end
  
  // How do we XOR the bits from our taps to generate the final feedback bit.
  // We can simply go over all bits and either XOR them or XOR a zero, XOR-ing a zero doesn't affect the output, its like multiplying by one.
  // we will chain each bit with the value of the previous bit's feedback XOR-ed either with it or with a zero if it is not a tap. 
  genvar i;
  generate  //  "generate" repetitive verilog code using loops instead.
    for(i=0; i < NUM_BITS; i = i+1) begin: lf   // So we loop over all the bits storing the current index inside i, we also name this loop lf (linear feedback) so that we will have a reference to access any wires or registers defined inside.
      wire feedback; // In each iteration of the loop we create a feedback wire and we connect it to one of two things. 
      if(i==0) // If we are on the first bit, there is no previous bit, so we simply take the current bit (sr[i]) AND-ed together with the same bit from the TAP parameter.
        assign feedback = sr[i] & TAPS[i]; // What this is doing is either evaluating to the value of current bit sr[i] if the TAP bit is 1, or making these two evaluate to zero if the TAP is not part of the XOR equation. By making it zero it won't affect the XOR operation.
      else
        assign feedback = lf[i-1].feedback ^ (sr[i] & TAPS[i]); // For all the other bits we take the previous feedback and XOR it with the same AND equation to either make it a zero if it is not part of our XOR equation, or return the value of sr[i].
    end
  endgenerate 
  assign finalFeedback = lf[NUM_BITS-1].feedback; // Take the output of the (last) XOR-ing. Connect the feedback from the final iteration to the wire we created finalFeedback: 
  // With that we now have a fully working LFSR of any size and any tap configuration.
endmodule