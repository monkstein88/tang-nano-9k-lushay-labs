module ROMBottom(input wire clk, input wire [10:0] addr, output reg [2:0] data = 0);

    always @(*) begin
        case (addr)
            11'b00000000000: data <= 3'b110;
            11'b00000000001: data <= 3'b110;
            11'b00000000010: data <= 3'b110;
            11'b00000000011: data <= 3'b110;
            11'b00000000100: data <= 3'b110;
            11'b00000000101: data <= 3'b110;
            11'b00000000110: data <= 3'b110;
            11'b00000000111: data <= 3'b110;
            11'b00000001000: data <= 3'b010;
            11'b00000001001: data <= 3'b110;
            11'b00000001010: data <= 3'b010;
            11'b00000001011: data <= 3'b011;
            11'b00000001100: data <= 3'b010;
            11'b00000001101: data <= 3'b010;
            11'b00000001110: data <= 3'b010;
            11'b00000001111: data <= 3'b011;
            11'b00000010000: data <= 3'b011;
            11'b00000010001: data <= 3'b011;
            11'b00000010010: data <= 3'b011;
            11'b00000010011: data <= 3'b010;
            11'b00000010100: data <= 3'b110;
            11'b00000010101: data <= 3'b110;
            11'b00000010110: data <= 3'b011;
            11'b00000010111: data <= 3'b011;
            11'b00000011000: data <= 3'b001;
            11'b00000011001: data <= 3'b001;
            11'b00000011010: data <= 3'b001;
            11'b00000011011: data <= 3'b001;
            11'b00000011100: data <= 3'b011;
            11'b00000011101: data <= 3'b011;
            11'b00000011110: data <= 3'b011;
            11'b00000011111: data <= 3'b011;
            11'b00000100000: data <= 3'b011;
            11'b00000100001: data <= 3'b011;
            11'b00000100010: data <= 3'b001;
            11'b00000100011: data <= 3'b001;
            11'b00000100100: data <= 3'b001;
            11'b00000100101: data <= 3'b001;
            11'b00000100110: data <= 3'b001;
            11'b00000100111: data <= 3'b011;
            11'b00000101000: data <= 3'b011;
            11'b00000101001: data <= 3'b010;
            11'b00000101010: data <= 3'b110;
            11'b00000101011: data <= 3'b010;
            11'b00000101100: data <= 3'b010;
            11'b00000101101: data <= 3'b011;
            11'b00000101110: data <= 3'b011;
            11'b00000101111: data <= 3'b011;
            11'b00000110000: data <= 3'b010;
            11'b00000110001: data <= 3'b010;
            11'b00000110010: data <= 3'b010;
            11'b00000110011: data <= 3'b011;
            11'b00000110100: data <= 3'b010;
            11'b00000110101: data <= 3'b110;
            11'b00000110110: data <= 3'b010;
            11'b00000110111: data <= 3'b110;
            11'b00000111000: data <= 3'b110;
            11'b00000111001: data <= 3'b110;
            11'b00000111010: data <= 3'b110;
            11'b00000111011: data <= 3'b110;
            11'b00000111100: data <= 3'b110;
            11'b00000111101: data <= 3'b110;
            11'b00000111110: data <= 3'b110;
            11'b00000111111: data <= 3'b110;
            11'b00001000000: data <= 3'b110;
            11'b00001000001: data <= 3'b110;
            11'b00001000010: data <= 3'b110;
            11'b00001000011: data <= 3'b110;
            11'b00001000100: data <= 3'b110;
            11'b00001000101: data <= 3'b110;
            11'b00001000110: data <= 3'b110;
            11'b00001000111: data <= 3'b110;
            11'b00001001000: data <= 3'b110;
            11'b00001001001: data <= 3'b110;
            11'b00001001010: data <= 3'b110;
            11'b00001001011: data <= 3'b010;
            11'b00001001100: data <= 3'b011;
            11'b00001001101: data <= 3'b011;
            11'b00001001110: data <= 3'b011;
            11'b00001001111: data <= 3'b011;
            11'b00001010000: data <= 3'b011;
            11'b00001010001: data <= 3'b011;
            11'b00001010010: data <= 3'b011;
            11'b00001010011: data <= 3'b011;
            11'b00001010100: data <= 3'b010;
            11'b00001010101: data <= 3'b010;
            11'b00001010110: data <= 3'b010;
            11'b00001010111: data <= 3'b011;
            11'b00001011000: data <= 3'b011;
            11'b00001011001: data <= 3'b001;
            11'b00001011010: data <= 3'b011;
            11'b00001011011: data <= 3'b011;
            11'b00001011100: data <= 3'b011;
            11'b00001011101: data <= 3'b011;
            11'b00001011110: data <= 3'b001;
            11'b00001011111: data <= 3'b001;
            11'b00001100000: data <= 3'b011;
            11'b00001100001: data <= 3'b011;
            11'b00001100010: data <= 3'b011;
            11'b00001100011: data <= 3'b011;
            11'b00001100100: data <= 3'b011;
            11'b00001100101: data <= 3'b001;
            11'b00001100110: data <= 3'b001;
            11'b00001100111: data <= 3'b011;
            11'b00001101000: data <= 3'b011;
            11'b00001101001: data <= 3'b010;
            11'b00001101010: data <= 3'b010;
            11'b00001101011: data <= 3'b011;
            11'b00001101100: data <= 3'b011;
            11'b00001101101: data <= 3'b011;
            11'b00001101110: data <= 3'b011;
            11'b00001101111: data <= 3'b011;
            11'b00001110000: data <= 3'b011;
            11'b00001110001: data <= 3'b011;
            11'b00001110010: data <= 3'b011;
            11'b00001110011: data <= 3'b010;
            11'b00001110100: data <= 3'b110;
            11'b00001110101: data <= 3'b110;
            11'b00001110110: data <= 3'b110;
            11'b00001110111: data <= 3'b110;
            11'b00001111000: data <= 3'b110;
            11'b00001111001: data <= 3'b110;
            11'b00001111010: data <= 3'b110;
            11'b00001111011: data <= 3'b110;
            11'b00001111100: data <= 3'b110;
            11'b00001111101: data <= 3'b110;
            11'b00001111110: data <= 3'b110;
            11'b00001111111: data <= 3'b110;
            11'b00010000000: data <= 3'b110;
            11'b00010000001: data <= 3'b110;
            11'b00010000010: data <= 3'b110;
            11'b00010000011: data <= 3'b110;
            11'b00010000100: data <= 3'b110;
            11'b00010000101: data <= 3'b110;
            11'b00010000110: data <= 3'b110;
            11'b00010000111: data <= 3'b110;
            11'b00010001000: data <= 3'b110;
            11'b00010001001: data <= 3'b110;
            11'b00010001010: data <= 3'b110;
            11'b00010001011: data <= 3'b110;
            11'b00010001100: data <= 3'b110;
            11'b00010001101: data <= 3'b010;
            11'b00010001110: data <= 3'b011;
            11'b00010001111: data <= 3'b011;
            11'b00010010000: data <= 3'b011;
            11'b00010010001: data <= 3'b011;
            11'b00010010010: data <= 3'b011;
            11'b00010010011: data <= 3'b011;
            11'b00010010100: data <= 3'b011;
            11'b00010010101: data <= 3'b011;
            11'b00010010110: data <= 3'b011;
            11'b00010010111: data <= 3'b011;
            11'b00010011000: data <= 3'b001;
            11'b00010011001: data <= 3'b001;
            11'b00010011010: data <= 3'b001;
            11'b00010011011: data <= 3'b001;
            11'b00010011100: data <= 3'b011;
            11'b00010011101: data <= 3'b011;
            11'b00010011110: data <= 3'b011;
            11'b00010011111: data <= 3'b001;
            11'b00010100000: data <= 3'b011;
            11'b00010100001: data <= 3'b011;
            11'b00010100010: data <= 3'b011;
            11'b00010100011: data <= 3'b011;
            11'b00010100100: data <= 3'b011;
            11'b00010100101: data <= 3'b001;
            11'b00010100110: data <= 3'b001;
            11'b00010100111: data <= 3'b011;
            11'b00010101000: data <= 3'b011;
            11'b00010101001: data <= 3'b011;
            11'b00010101010: data <= 3'b011;
            11'b00010101011: data <= 3'b011;
            11'b00010101100: data <= 3'b011;
            11'b00010101101: data <= 3'b011;
            11'b00010101110: data <= 3'b011;
            11'b00010101111: data <= 3'b011;
            11'b00010110000: data <= 3'b011;
            11'b00010110001: data <= 3'b010;
            11'b00010110010: data <= 3'b110;
            11'b00010110011: data <= 3'b110;
            11'b00010110100: data <= 3'b110;
            11'b00010110101: data <= 3'b110;
            11'b00010110110: data <= 3'b110;
            11'b00010110111: data <= 3'b110;
            11'b00010111000: data <= 3'b110;
            11'b00010111001: data <= 3'b110;
            11'b00010111010: data <= 3'b110;
            11'b00010111011: data <= 3'b110;
            11'b00010111100: data <= 3'b110;
            11'b00010111101: data <= 3'b110;
            11'b00010111110: data <= 3'b110;
            11'b00010111111: data <= 3'b110;
            11'b00011000000: data <= 3'b110;
            11'b00011000001: data <= 3'b110;
            11'b00011000010: data <= 3'b110;
            11'b00011000011: data <= 3'b110;
            11'b00011000100: data <= 3'b110;
            11'b00011000101: data <= 3'b110;
            11'b00011000110: data <= 3'b110;
            11'b00011000111: data <= 3'b110;
            11'b00011001000: data <= 3'b110;
            11'b00011001001: data <= 3'b110;
            11'b00011001010: data <= 3'b110;
            11'b00011001011: data <= 3'b110;
            11'b00011001100: data <= 3'b110;
            11'b00011001101: data <= 3'b010;
            11'b00011001110: data <= 3'b011;
            11'b00011001111: data <= 3'b011;
            11'b00011010000: data <= 3'b011;
            11'b00011010001: data <= 3'b010;
            11'b00011010010: data <= 3'b010;
            11'b00011010011: data <= 3'b011;
            11'b00011010100: data <= 3'b011;
            11'b00011010101: data <= 3'b011;
            11'b00011010110: data <= 3'b011;
            11'b00011010111: data <= 3'b011;
            11'b00011011000: data <= 3'b011;
            11'b00011011001: data <= 3'b001;
            11'b00011011010: data <= 3'b001;
            11'b00011011011: data <= 3'b011;
            11'b00011011100: data <= 3'b001;
            11'b00011011101: data <= 3'b011;
            11'b00011011110: data <= 3'b011;
            11'b00011011111: data <= 3'b001;
            11'b00011100000: data <= 3'b001;
            11'b00011100001: data <= 3'b001;
            11'b00011100010: data <= 3'b001;
            11'b00011100011: data <= 3'b011;
            11'b00011100100: data <= 3'b001;
            11'b00011100101: data <= 3'b001;
            11'b00011100110: data <= 3'b011;
            11'b00011100111: data <= 3'b010;
            11'b00011101000: data <= 3'b011;
            11'b00011101001: data <= 3'b011;
            11'b00011101010: data <= 3'b011;
            11'b00011101011: data <= 3'b011;
            11'b00011101100: data <= 3'b011;
            11'b00011101101: data <= 3'b010;
            11'b00011101110: data <= 3'b011;
            11'b00011101111: data <= 3'b011;
            11'b00011110000: data <= 3'b011;
            11'b00011110001: data <= 3'b010;
            11'b00011110010: data <= 3'b110;
            11'b00011110011: data <= 3'b110;
            11'b00011110100: data <= 3'b110;
            11'b00011110101: data <= 3'b110;
            11'b00011110110: data <= 3'b110;
            11'b00011110111: data <= 3'b110;
            11'b00011111000: data <= 3'b110;
            11'b00011111001: data <= 3'b110;
            11'b00011111010: data <= 3'b110;
            11'b00011111011: data <= 3'b110;
            11'b00011111100: data <= 3'b110;
            11'b00011111101: data <= 3'b110;
            11'b00011111110: data <= 3'b110;
            11'b00011111111: data <= 3'b110;
            11'b00100000000: data <= 3'b110;
            11'b00100000001: data <= 3'b110;
            11'b00100000010: data <= 3'b110;
            11'b00100000011: data <= 3'b110;
            11'b00100000100: data <= 3'b110;
            11'b00100000101: data <= 3'b110;
            11'b00100000110: data <= 3'b110;
            11'b00100000111: data <= 3'b110;
            11'b00100001000: data <= 3'b110;
            11'b00100001001: data <= 3'b110;
            11'b00100001010: data <= 3'b110;
            11'b00100001011: data <= 3'b010;
            11'b00100001100: data <= 3'b011;
            11'b00100001101: data <= 3'b011;
            11'b00100001110: data <= 3'b011;
            11'b00100001111: data <= 3'b011;
            11'b00100010000: data <= 3'b011;
            11'b00100010001: data <= 3'b110;
            11'b00100010010: data <= 3'b110;
            11'b00100010011: data <= 3'b011;
            11'b00100010100: data <= 3'b011;
            11'b00100010101: data <= 3'b011;
            11'b00100010110: data <= 3'b011;
            11'b00100010111: data <= 3'b010;
            11'b00100011000: data <= 3'b011;
            11'b00100011001: data <= 3'b001;
            11'b00100011010: data <= 3'b011;
            11'b00100011011: data <= 3'b011;
            11'b00100011100: data <= 3'b011;
            11'b00100011101: data <= 3'b011;
            11'b00100011110: data <= 3'b001;
            11'b00100011111: data <= 3'b001;
            11'b00100100000: data <= 3'b001;
            11'b00100100001: data <= 3'b011;
            11'b00100100010: data <= 3'b011;
            11'b00100100011: data <= 3'b011;
            11'b00100100100: data <= 3'b011;
            11'b00100100101: data <= 3'b001;
            11'b00100100110: data <= 3'b011;
            11'b00100100111: data <= 3'b010;
            11'b00100101000: data <= 3'b011;
            11'b00100101001: data <= 3'b011;
            11'b00100101010: data <= 3'b011;
            11'b00100101011: data <= 3'b011;
            11'b00100101100: data <= 3'b010;
            11'b00100101101: data <= 3'b110;
            11'b00100101110: data <= 3'b010;
            11'b00100101111: data <= 3'b011;
            11'b00100110000: data <= 3'b011;
            11'b00100110001: data <= 3'b011;
            11'b00100110010: data <= 3'b011;
            11'b00100110011: data <= 3'b011;
            11'b00100110100: data <= 3'b010;
            11'b00100110101: data <= 3'b110;
            11'b00100110110: data <= 3'b110;
            11'b00100110111: data <= 3'b110;
            11'b00100111000: data <= 3'b110;
            11'b00100111001: data <= 3'b110;
            11'b00100111010: data <= 3'b110;
            11'b00100111011: data <= 3'b110;
            11'b00100111100: data <= 3'b110;
            11'b00100111101: data <= 3'b110;
            11'b00100111110: data <= 3'b110;
            11'b00100111111: data <= 3'b110;
            11'b00101000000: data <= 3'b110;
            11'b00101000001: data <= 3'b110;
            11'b00101000010: data <= 3'b110;
            11'b00101000011: data <= 3'b110;
            11'b00101000100: data <= 3'b110;
            11'b00101000101: data <= 3'b110;
            11'b00101000110: data <= 3'b110;
            11'b00101000111: data <= 3'b110;
            11'b00101001000: data <= 3'b110;
            11'b00101001001: data <= 3'b010;
            11'b00101001010: data <= 3'b011;
            11'b00101001011: data <= 3'b011;
            11'b00101001100: data <= 3'b011;
            11'b00101001101: data <= 3'b011;
            11'b00101001110: data <= 3'b011;
            11'b00101001111: data <= 3'b011;
            11'b00101010000: data <= 3'b010;
            11'b00101010001: data <= 3'b110;
            11'b00101010010: data <= 3'b010;
            11'b00101010011: data <= 3'b011;
            11'b00101010100: data <= 3'b011;
            11'b00101010101: data <= 3'b011;
            11'b00101010110: data <= 3'b010;
            11'b00101010111: data <= 3'b110;
            11'b00101011000: data <= 3'b010;
            11'b00101011001: data <= 3'b011;
            11'b00101011010: data <= 3'b001;
            11'b00101011011: data <= 3'b011;
            11'b00101011100: data <= 3'b011;
            11'b00101011101: data <= 3'b001;
            11'b00101011110: data <= 3'b001;
            11'b00101011111: data <= 3'b001;
            11'b00101100000: data <= 3'b001;
            11'b00101100001: data <= 3'b001;
            11'b00101100010: data <= 3'b011;
            11'b00101100011: data <= 3'b001;
            11'b00101100100: data <= 3'b001;
            11'b00101100101: data <= 3'b001;
            11'b00101100110: data <= 3'b010;
            11'b00101100111: data <= 3'b110;
            11'b00101101000: data <= 3'b010;
            11'b00101101001: data <= 3'b011;
            11'b00101101010: data <= 3'b011;
            11'b00101101011: data <= 3'b011;
            11'b00101101100: data <= 3'b010;
            11'b00101101101: data <= 3'b110;
            11'b00101101110: data <= 3'b010;
            11'b00101101111: data <= 3'b011;
            11'b00101110000: data <= 3'b011;
            11'b00101110001: data <= 3'b011;
            11'b00101110010: data <= 3'b011;
            11'b00101110011: data <= 3'b011;
            11'b00101110100: data <= 3'b011;
            11'b00101110101: data <= 3'b010;
            11'b00101110110: data <= 3'b110;
            11'b00101110111: data <= 3'b110;
            11'b00101111000: data <= 3'b110;
            11'b00101111001: data <= 3'b110;
            11'b00101111010: data <= 3'b110;
            11'b00101111011: data <= 3'b110;
            11'b00101111100: data <= 3'b110;
            11'b00101111101: data <= 3'b110;
            11'b00101111110: data <= 3'b110;
            11'b00101111111: data <= 3'b110;
            11'b00110000000: data <= 3'b110;
            11'b00110000001: data <= 3'b110;
            11'b00110000010: data <= 3'b110;
            11'b00110000011: data <= 3'b110;
            11'b00110000100: data <= 3'b110;
            11'b00110000101: data <= 3'b110;
            11'b00110000110: data <= 3'b010;
            11'b00110000111: data <= 3'b010;
            11'b00110001000: data <= 3'b110;
            11'b00110001001: data <= 3'b010;
            11'b00110001010: data <= 3'b011;
            11'b00110001011: data <= 3'b011;
            11'b00110001100: data <= 3'b011;
            11'b00110001101: data <= 3'b010;
            11'b00110001110: data <= 3'b010;
            11'b00110001111: data <= 3'b010;
            11'b00110010000: data <= 3'b010;
            11'b00110010001: data <= 3'b010;
            11'b00110010010: data <= 3'b010;
            11'b00110010011: data <= 3'b011;
            11'b00110010100: data <= 3'b011;
            11'b00110010101: data <= 3'b011;
            11'b00110010110: data <= 3'b011;
            11'b00110010111: data <= 3'b010;
            11'b00110011000: data <= 3'b010;
            11'b00110011001: data <= 3'b011;
            11'b00110011010: data <= 3'b010;
            11'b00110011011: data <= 3'b000;
            11'b00110011100: data <= 3'b001;
            11'b00110011101: data <= 3'b001;
            11'b00110011110: data <= 3'b001;
            11'b00110011111: data <= 3'b001;
            11'b00110100000: data <= 3'b001;
            11'b00110100001: data <= 3'b001;
            11'b00110100010: data <= 3'b001;
            11'b00110100011: data <= 3'b000;
            11'b00110100100: data <= 3'b010;
            11'b00110100101: data <= 3'b011;
            11'b00110100110: data <= 3'b010;
            11'b00110100111: data <= 3'b110;
            11'b00110101000: data <= 3'b010;
            11'b00110101001: data <= 3'b011;
            11'b00110101010: data <= 3'b011;
            11'b00110101011: data <= 3'b011;
            11'b00110101100: data <= 3'b010;
            11'b00110101101: data <= 3'b010;
            11'b00110101110: data <= 3'b010;
            11'b00110101111: data <= 3'b010;
            11'b00110110000: data <= 3'b010;
            11'b00110110001: data <= 3'b010;
            11'b00110110010: data <= 3'b011;
            11'b00110110011: data <= 3'b011;
            11'b00110110100: data <= 3'b011;
            11'b00110110101: data <= 3'b011;
            11'b00110110110: data <= 3'b110;
            11'b00110110111: data <= 3'b010;
            11'b00110111000: data <= 3'b010;
            11'b00110111001: data <= 3'b110;
            11'b00110111010: data <= 3'b110;
            11'b00110111011: data <= 3'b110;
            11'b00110111100: data <= 3'b110;
            11'b00110111101: data <= 3'b110;
            11'b00110111110: data <= 3'b110;
            11'b00110111111: data <= 3'b110;
            11'b00111000000: data <= 3'b110;
            11'b00111000001: data <= 3'b110;
            11'b00111000010: data <= 3'b110;
            11'b00111000011: data <= 3'b110;
            11'b00111000100: data <= 3'b110;
            11'b00111000101: data <= 3'b110;
            11'b00111000110: data <= 3'b010;
            11'b00111000111: data <= 3'b010;
            11'b00111001000: data <= 3'b010;
            11'b00111001001: data <= 3'b010;
            11'b00111001010: data <= 3'b010;
            11'b00111001011: data <= 3'b011;
            11'b00111001100: data <= 3'b011;
            11'b00111001101: data <= 3'b110;
            11'b00111001110: data <= 3'b010;
            11'b00111001111: data <= 3'b010;
            11'b00111010000: data <= 3'b010;
            11'b00111010001: data <= 3'b010;
            11'b00111010010: data <= 3'b010;
            11'b00111010011: data <= 3'b010;
            11'b00111010100: data <= 3'b010;
            11'b00111010101: data <= 3'b011;
            11'b00111010110: data <= 3'b011;
            11'b00111010111: data <= 3'b011;
            11'b00111011000: data <= 3'b011;
            11'b00111011001: data <= 3'b011;
            11'b00111011010: data <= 3'b110;
            11'b00111011011: data <= 3'b110;
            11'b00111011100: data <= 3'b010;
            11'b00111011101: data <= 3'b001;
            11'b00111011110: data <= 3'b001;
            11'b00111011111: data <= 3'b001;
            11'b00111100000: data <= 3'b001;
            11'b00111100001: data <= 3'b001;
            11'b00111100010: data <= 3'b010;
            11'b00111100011: data <= 3'b110;
            11'b00111100100: data <= 3'b010;
            11'b00111100101: data <= 3'b010;
            11'b00111100110: data <= 3'b011;
            11'b00111100111: data <= 3'b011;
            11'b00111101000: data <= 3'b011;
            11'b00111101001: data <= 3'b011;
            11'b00111101010: data <= 3'b010;
            11'b00111101011: data <= 3'b010;
            11'b00111101100: data <= 3'b010;
            11'b00111101101: data <= 3'b010;
            11'b00111101110: data <= 3'b010;
            11'b00111101111: data <= 3'b010;
            11'b00111110000: data <= 3'b010;
            11'b00111110001: data <= 3'b110;
            11'b00111110010: data <= 3'b011;
            11'b00111110011: data <= 3'b011;
            11'b00111110100: data <= 3'b010;
            11'b00111110101: data <= 3'b010;
            11'b00111110110: data <= 3'b010;
            11'b00111110111: data <= 3'b010;
            11'b00111111000: data <= 3'b010;
            11'b00111111001: data <= 3'b010;
            11'b00111111010: data <= 3'b110;
            11'b00111111011: data <= 3'b110;
            11'b00111111100: data <= 3'b110;
            11'b00111111101: data <= 3'b110;
            11'b00111111110: data <= 3'b110;
            11'b00111111111: data <= 3'b110;
            11'b01000000000: data <= 3'b010;
            11'b01000000001: data <= 3'b010;
            11'b01000000010: data <= 3'b010;
            11'b01000000011: data <= 3'b010;
            11'b01000000100: data <= 3'b010;
            11'b01000000101: data <= 3'b010;
            11'b01000000110: data <= 3'b010;
            11'b01000000111: data <= 3'b010;
            11'b01000001000: data <= 3'b010;
            11'b01000001001: data <= 3'b010;
            11'b01000001010: data <= 3'b010;
            11'b01000001011: data <= 3'b011;
            11'b01000001100: data <= 3'b011;
            11'b01000001101: data <= 3'b011;
            11'b01000001110: data <= 3'b011;
            11'b01000001111: data <= 3'b010;
            11'b01000010000: data <= 3'b010;
            11'b01000010001: data <= 3'b010;
            11'b01000010010: data <= 3'b010;
            11'b01000010011: data <= 3'b010;
            11'b01000010100: data <= 3'b110;
            11'b01000010101: data <= 3'b010;
            11'b01000010110: data <= 3'b011;
            11'b01000010111: data <= 3'b011;
            11'b01000011000: data <= 3'b011;
            11'b01000011001: data <= 3'b010;
            11'b01000011010: data <= 3'b010;
            11'b01000011011: data <= 3'b010;
            11'b01000011100: data <= 3'b010;
            11'b01000011101: data <= 3'b010;
            11'b01000011110: data <= 3'b011;
            11'b01000011111: data <= 3'b011;
            11'b01000100000: data <= 3'b011;
            11'b01000100001: data <= 3'b010;
            11'b01000100010: data <= 3'b010;
            11'b01000100011: data <= 3'b010;
            11'b01000100100: data <= 3'b010;
            11'b01000100101: data <= 3'b010;
            11'b01000100110: data <= 3'b011;
            11'b01000100111: data <= 3'b011;
            11'b01000101000: data <= 3'b011;
            11'b01000101001: data <= 3'b010;
            11'b01000101010: data <= 3'b110;
            11'b01000101011: data <= 3'b010;
            11'b01000101100: data <= 3'b010;
            11'b01000101101: data <= 3'b010;
            11'b01000101110: data <= 3'b010;
            11'b01000101111: data <= 3'b110;
            11'b01000110000: data <= 3'b011;
            11'b01000110001: data <= 3'b011;
            11'b01000110010: data <= 3'b011;
            11'b01000110011: data <= 3'b011;
            11'b01000110100: data <= 3'b010;
            11'b01000110101: data <= 3'b010;
            11'b01000110110: data <= 3'b010;
            11'b01000110111: data <= 3'b010;
            11'b01000111000: data <= 3'b010;
            11'b01000111001: data <= 3'b010;
            11'b01000111010: data <= 3'b010;
            11'b01000111011: data <= 3'b010;
            11'b01000111100: data <= 3'b010;
            11'b01000111101: data <= 3'b010;
            11'b01000111110: data <= 3'b010;
            11'b01000111111: data <= 3'b010;
            11'b01001000000: data <= 3'b110;
            11'b01001000001: data <= 3'b110;
            11'b01001000010: data <= 3'b110;
            11'b01001000011: data <= 3'b110;
            11'b01001000100: data <= 3'b110;
            11'b01001000101: data <= 3'b110;
            11'b01001000110: data <= 3'b110;
            11'b01001000111: data <= 3'b010;
            11'b01001001000: data <= 3'b010;
            11'b01001001001: data <= 3'b110;
            11'b01001001010: data <= 3'b010;
            11'b01001001011: data <= 3'b011;
            11'b01001001100: data <= 3'b011;
            11'b01001001101: data <= 3'b011;
            11'b01001001110: data <= 3'b011;
            11'b01001001111: data <= 3'b010;
            11'b01001010000: data <= 3'b010;
            11'b01001010001: data <= 3'b010;
            11'b01001010010: data <= 3'b010;
            11'b01001010011: data <= 3'b010;
            11'b01001010100: data <= 3'b010;
            11'b01001010101: data <= 3'b011;
            11'b01001010110: data <= 3'b011;
            11'b01001010111: data <= 3'b010;
            11'b01001011000: data <= 3'b010;
            11'b01001011001: data <= 3'b010;
            11'b01001011010: data <= 3'b010;
            11'b01001011011: data <= 3'b010;
            11'b01001011100: data <= 3'b010;
            11'b01001011101: data <= 3'b010;
            11'b01001011110: data <= 3'b010;
            11'b01001011111: data <= 3'b010;
            11'b01001100000: data <= 3'b010;
            11'b01001100001: data <= 3'b010;
            11'b01001100010: data <= 3'b010;
            11'b01001100011: data <= 3'b010;
            11'b01001100100: data <= 3'b010;
            11'b01001100101: data <= 3'b010;
            11'b01001100110: data <= 3'b010;
            11'b01001100111: data <= 3'b010;
            11'b01001101000: data <= 3'b011;
            11'b01001101001: data <= 3'b011;
            11'b01001101010: data <= 3'b010;
            11'b01001101011: data <= 3'b010;
            11'b01001101100: data <= 3'b010;
            11'b01001101101: data <= 3'b010;
            11'b01001101110: data <= 3'b010;
            11'b01001101111: data <= 3'b010;
            11'b01001110000: data <= 3'b010;
            11'b01001110001: data <= 3'b011;
            11'b01001110010: data <= 3'b011;
            11'b01001110011: data <= 3'b011;
            11'b01001110100: data <= 3'b010;
            11'b01001110101: data <= 3'b110;
            11'b01001110110: data <= 3'b010;
            11'b01001110111: data <= 3'b010;
            11'b01001111000: data <= 3'b110;
            11'b01001111001: data <= 3'b110;
            11'b01001111010: data <= 3'b110;
            11'b01001111011: data <= 3'b110;
            11'b01001111100: data <= 3'b110;
            11'b01001111101: data <= 3'b110;
            11'b01001111110: data <= 3'b110;
            11'b01001111111: data <= 3'b110;
            11'b01010000000: data <= 3'b010;
            11'b01010000001: data <= 3'b010;
            11'b01010000010: data <= 3'b010;
            11'b01010000011: data <= 3'b010;
            11'b01010000100: data <= 3'b010;
            11'b01010000101: data <= 3'b010;
            11'b01010000110: data <= 3'b010;
            11'b01010000111: data <= 3'b010;
            11'b01010001000: data <= 3'b010;
            11'b01010001001: data <= 3'b010;
            11'b01010001010: data <= 3'b011;
            11'b01010001011: data <= 3'b010;
            11'b01010001100: data <= 3'b010;
            11'b01010001101: data <= 3'b010;
            11'b01010001110: data <= 3'b011;
            11'b01010001111: data <= 3'b011;
            11'b01010010000: data <= 3'b010;
            11'b01010010001: data <= 3'b110;
            11'b01010010010: data <= 3'b111;
            11'b01010010011: data <= 3'b110;
            11'b01010010100: data <= 3'b000;
            11'b01010010101: data <= 3'b011;
            11'b01010010110: data <= 3'b011;
            11'b01010010111: data <= 3'b000;
            11'b01010011000: data <= 3'b010;
            11'b01010011001: data <= 3'b010;
            11'b01010011010: data <= 3'b010;
            11'b01010011011: data <= 3'b010;
            11'b01010011100: data <= 3'b010;
            11'b01010011101: data <= 3'b110;
            11'b01010011110: data <= 3'b010;
            11'b01010011111: data <= 3'b010;
            11'b01010100000: data <= 3'b010;
            11'b01010100001: data <= 3'b110;
            11'b01010100010: data <= 3'b010;
            11'b01010100011: data <= 3'b010;
            11'b01010100100: data <= 3'b010;
            11'b01010100101: data <= 3'b010;
            11'b01010100110: data <= 3'b010;
            11'b01010100111: data <= 3'b000;
            11'b01010101000: data <= 3'b010;
            11'b01010101001: data <= 3'b011;
            11'b01010101010: data <= 3'b000;
            11'b01010101011: data <= 3'b110;
            11'b01010101100: data <= 3'b111;
            11'b01010101101: data <= 3'b110;
            11'b01010101110: data <= 3'b000;
            11'b01010101111: data <= 3'b011;
            11'b01010110000: data <= 3'b011;
            11'b01010110001: data <= 3'b010;
            11'b01010110010: data <= 3'b010;
            11'b01010110011: data <= 3'b010;
            11'b01010110100: data <= 3'b011;
            11'b01010110101: data <= 3'b010;
            11'b01010110110: data <= 3'b010;
            11'b01010110111: data <= 3'b010;
            11'b01010111000: data <= 3'b010;
            11'b01010111001: data <= 3'b010;
            11'b01010111010: data <= 3'b010;
            11'b01010111011: data <= 3'b010;
            11'b01010111100: data <= 3'b010;
            11'b01010111101: data <= 3'b010;
            11'b01010111110: data <= 3'b010;
            11'b01010111111: data <= 3'b010;
            11'b01011000000: data <= 3'b001;
            11'b01011000001: data <= 3'b001;
            11'b01011000010: data <= 3'b001;
            11'b01011000011: data <= 3'b001;
            11'b01011000100: data <= 3'b001;
            11'b01011000101: data <= 3'b001;
            11'b01011000110: data <= 3'b001;
            11'b01011000111: data <= 3'b010;
            11'b01011001000: data <= 3'b010;
            11'b01011001001: data <= 3'b011;
            11'b01011001010: data <= 3'b011;
            11'b01011001011: data <= 3'b010;
            11'b01011001100: data <= 3'b010;
            11'b01011001101: data <= 3'b010;
            11'b01011001110: data <= 3'b010;
            11'b01011001111: data <= 3'b011;
            11'b01011010000: data <= 3'b001;
            11'b01011010001: data <= 3'b111;
            11'b01011010010: data <= 3'b111;
            11'b01011010011: data <= 3'b111;
            11'b01011010100: data <= 3'b011;
            11'b01011010101: data <= 3'b001;
            11'b01011010110: data <= 3'b001;
            11'b01011010111: data <= 3'b110;
            11'b01011011000: data <= 3'b010;
            11'b01011011001: data <= 3'b010;
            11'b01011011010: data <= 3'b010;
            11'b01011011011: data <= 3'b010;
            11'b01011011100: data <= 3'b010;
            11'b01011011101: data <= 3'b000;
            11'b01011011110: data <= 3'b010;
            11'b01011011111: data <= 3'b010;
            11'b01011100000: data <= 3'b010;
            11'b01011100001: data <= 3'b000;
            11'b01011100010: data <= 3'b010;
            11'b01011100011: data <= 3'b010;
            11'b01011100100: data <= 3'b010;
            11'b01011100101: data <= 3'b010;
            11'b01011100110: data <= 3'b010;
            11'b01011100111: data <= 3'b110;
            11'b01011101000: data <= 3'b001;
            11'b01011101001: data <= 3'b001;
            11'b01011101010: data <= 3'b011;
            11'b01011101011: data <= 3'b111;
            11'b01011101100: data <= 3'b111;
            11'b01011101101: data <= 3'b001;
            11'b01011101110: data <= 3'b001;
            11'b01011101111: data <= 3'b011;
            11'b01011110000: data <= 3'b010;
            11'b01011110001: data <= 3'b010;
            11'b01011110010: data <= 3'b010;
            11'b01011110011: data <= 3'b010;
            11'b01011110100: data <= 3'b011;
            11'b01011110101: data <= 3'b011;
            11'b01011110110: data <= 3'b010;
            11'b01011110111: data <= 3'b010;
            11'b01011111000: data <= 3'b001;
            11'b01011111001: data <= 3'b001;
            11'b01011111010: data <= 3'b001;
            11'b01011111011: data <= 3'b001;
            11'b01011111100: data <= 3'b001;
            11'b01011111101: data <= 3'b001;
            11'b01011111110: data <= 3'b001;
            11'b01011111111: data <= 3'b001;
            11'b01100000000: data <= 3'b001;
            11'b01100000001: data <= 3'b001;
            11'b01100000010: data <= 3'b001;
            11'b01100000011: data <= 3'b001;
            11'b01100000100: data <= 3'b001;
            11'b01100000101: data <= 3'b001;
            11'b01100000110: data <= 3'b001;
            11'b01100000111: data <= 3'b001;
            11'b01100001000: data <= 3'b000;
            11'b01100001001: data <= 3'b010;
            11'b01100001010: data <= 3'b010;
            11'b01100001011: data <= 3'b010;
            11'b01100001100: data <= 3'b010;
            11'b01100001101: data <= 3'b010;
            11'b01100001110: data <= 3'b010;
            11'b01100001111: data <= 3'b010;
            11'b01100010000: data <= 3'b010;
            11'b01100010001: data <= 3'b000;
            11'b01100010010: data <= 3'b001;
            11'b01100010011: data <= 3'b111;
            11'b01100010100: data <= 3'b111;
            11'b01100010101: data <= 3'b111;
            11'b01100010110: data <= 3'b001;
            11'b01100010111: data <= 3'b000;
            11'b01100011000: data <= 3'b000;
            11'b01100011001: data <= 3'b010;
            11'b01100011010: data <= 3'b010;
            11'b01100011011: data <= 3'b010;
            11'b01100011100: data <= 3'b000;
            11'b01100011101: data <= 3'b010;
            11'b01100011110: data <= 3'b010;
            11'b01100011111: data <= 3'b001;
            11'b01100100000: data <= 3'b010;
            11'b01100100001: data <= 3'b010;
            11'b01100100010: data <= 3'b000;
            11'b01100100011: data <= 3'b010;
            11'b01100100100: data <= 3'b010;
            11'b01100100101: data <= 3'b010;
            11'b01100100110: data <= 3'b000;
            11'b01100100111: data <= 3'b000;
            11'b01100101000: data <= 3'b001;
            11'b01100101001: data <= 3'b111;
            11'b01100101010: data <= 3'b111;
            11'b01100101011: data <= 3'b111;
            11'b01100101100: data <= 3'b001;
            11'b01100101101: data <= 3'b000;
            11'b01100101110: data <= 3'b110;
            11'b01100101111: data <= 3'b010;
            11'b01100110000: data <= 3'b010;
            11'b01100110001: data <= 3'b010;
            11'b01100110010: data <= 3'b010;
            11'b01100110011: data <= 3'b010;
            11'b01100110100: data <= 3'b010;
            11'b01100110101: data <= 3'b010;
            11'b01100110110: data <= 3'b000;
            11'b01100110111: data <= 3'b001;
            11'b01100111000: data <= 3'b001;
            11'b01100111001: data <= 3'b001;
            11'b01100111010: data <= 3'b001;
            11'b01100111011: data <= 3'b001;
            11'b01100111100: data <= 3'b001;
            11'b01100111101: data <= 3'b001;
            11'b01100111110: data <= 3'b001;
            11'b01100111111: data <= 3'b001;
            11'b01101000000: data <= 3'b001;
            11'b01101000001: data <= 3'b001;
            11'b01101000010: data <= 3'b001;
            11'b01101000011: data <= 3'b001;
            11'b01101000100: data <= 3'b001;
            11'b01101000101: data <= 3'b001;
            11'b01101000110: data <= 3'b001;
            11'b01101000111: data <= 3'b001;
            11'b01101001000: data <= 3'b001;
            11'b01101001001: data <= 3'b000;
            11'b01101001010: data <= 3'b110;
            11'b01101001011: data <= 3'b010;
            11'b01101001100: data <= 3'b010;
            11'b01101001101: data <= 3'b010;
            11'b01101001110: data <= 3'b010;
            11'b01101001111: data <= 3'b010;
            11'b01101010000: data <= 3'b110;
            11'b01101010001: data <= 3'b111;
            11'b01101010010: data <= 3'b000;
            11'b01101010011: data <= 3'b001;
            11'b01101010100: data <= 3'b111;
            11'b01101010101: data <= 3'b111;
            11'b01101010110: data <= 3'b111;
            11'b01101010111: data <= 3'b001;
            11'b01101011000: data <= 3'b001;
            11'b01101011001: data <= 3'b001;
            11'b01101011010: data <= 3'b001;
            11'b01101011011: data <= 3'b000;
            11'b01101011100: data <= 3'b010;
            11'b01101011101: data <= 3'b010;
            11'b01101011110: data <= 3'b001;
            11'b01101011111: data <= 3'b001;
            11'b01101100000: data <= 3'b001;
            11'b01101100001: data <= 3'b010;
            11'b01101100010: data <= 3'b110;
            11'b01101100011: data <= 3'b010;
            11'b01101100100: data <= 3'b001;
            11'b01101100101: data <= 3'b001;
            11'b01101100110: data <= 3'b001;
            11'b01101100111: data <= 3'b001;
            11'b01101101000: data <= 3'b111;
            11'b01101101001: data <= 3'b111;
            11'b01101101010: data <= 3'b111;
            11'b01101101011: data <= 3'b001;
            11'b01101101100: data <= 3'b001;
            11'b01101101101: data <= 3'b111;
            11'b01101101110: data <= 3'b110;
            11'b01101101111: data <= 3'b010;
            11'b01101110000: data <= 3'b010;
            11'b01101110001: data <= 3'b010;
            11'b01101110010: data <= 3'b010;
            11'b01101110011: data <= 3'b010;
            11'b01101110100: data <= 3'b110;
            11'b01101110101: data <= 3'b000;
            11'b01101110110: data <= 3'b001;
            11'b01101110111: data <= 3'b001;
            11'b01101111000: data <= 3'b001;
            11'b01101111001: data <= 3'b001;
            11'b01101111010: data <= 3'b001;
            11'b01101111011: data <= 3'b001;
            11'b01101111100: data <= 3'b001;
            11'b01101111101: data <= 3'b001;
            11'b01101111110: data <= 3'b001;
            11'b01101111111: data <= 3'b001;
            11'b01110000000: data <= 3'b001;
            11'b01110000001: data <= 3'b001;
            11'b01110000010: data <= 3'b001;
            11'b01110000011: data <= 3'b001;
            11'b01110000100: data <= 3'b001;
            11'b01110000101: data <= 3'b001;
            11'b01110000110: data <= 3'b001;
            11'b01110000111: data <= 3'b001;
            11'b01110001000: data <= 3'b001;
            11'b01110001001: data <= 3'b001;
            11'b01110001010: data <= 3'b000;
            11'b01110001011: data <= 3'b000;
            11'b01110001100: data <= 3'b001;
            11'b01110001101: data <= 3'b000;
            11'b01110001110: data <= 3'b110;
            11'b01110001111: data <= 3'b010;
            11'b01110010000: data <= 3'b110;
            11'b01110010001: data <= 3'b111;
            11'b01110010010: data <= 3'b111;
            11'b01110010011: data <= 3'b111;
            11'b01110010100: data <= 3'b111;
            11'b01110010101: data <= 3'b000;
            11'b01110010110: data <= 3'b111;
            11'b01110010111: data <= 3'b111;
            11'b01110011000: data <= 3'b111;
            11'b01110011001: data <= 3'b000;
            11'b01110011010: data <= 3'b000;
            11'b01110011011: data <= 3'b000;
            11'b01110011100: data <= 3'b000;
            11'b01110011101: data <= 3'b001;
            11'b01110011110: data <= 3'b001;
            11'b01110011111: data <= 3'b001;
            11'b01110100000: data <= 3'b001;
            11'b01110100001: data <= 3'b001;
            11'b01110100010: data <= 3'b001;
            11'b01110100011: data <= 3'b000;
            11'b01110100100: data <= 3'b001;
            11'b01110100101: data <= 3'b001;
            11'b01110100110: data <= 3'b111;
            11'b01110100111: data <= 3'b111;
            11'b01110101000: data <= 3'b111;
            11'b01110101001: data <= 3'b011;
            11'b01110101010: data <= 3'b111;
            11'b01110101011: data <= 3'b111;
            11'b01110101100: data <= 3'b111;
            11'b01110101101: data <= 3'b111;
            11'b01110101110: data <= 3'b110;
            11'b01110101111: data <= 3'b010;
            11'b01110110000: data <= 3'b110;
            11'b01110110001: data <= 3'b000;
            11'b01110110010: data <= 3'b001;
            11'b01110110011: data <= 3'b000;
            11'b01110110100: data <= 3'b000;
            11'b01110110101: data <= 3'b001;
            11'b01110110110: data <= 3'b001;
            11'b01110110111: data <= 3'b001;
            11'b01110111000: data <= 3'b001;
            11'b01110111001: data <= 3'b001;
            11'b01110111010: data <= 3'b001;
            11'b01110111011: data <= 3'b001;
            11'b01110111100: data <= 3'b001;
            11'b01110111101: data <= 3'b001;
            11'b01110111110: data <= 3'b001;
            11'b01110111111: data <= 3'b001;
            11'b01111000000: data <= 3'b001;
            11'b01111000001: data <= 3'b001;
            11'b01111000010: data <= 3'b001;
            11'b01111000011: data <= 3'b001;
            11'b01111000100: data <= 3'b001;
            11'b01111000101: data <= 3'b001;
            11'b01111000110: data <= 3'b001;
            11'b01111000111: data <= 3'b001;
            11'b01111001000: data <= 3'b001;
            11'b01111001001: data <= 3'b001;
            11'b01111001010: data <= 3'b001;
            11'b01111001011: data <= 3'b001;
            11'b01111001100: data <= 3'b001;
            11'b01111001101: data <= 3'b010;
            11'b01111001110: data <= 3'b110;
            11'b01111001111: data <= 3'b001;
            11'b01111010000: data <= 3'b001;
            11'b01111010001: data <= 3'b111;
            11'b01111010010: data <= 3'b111;
            11'b01111010011: data <= 3'b011;
            11'b01111010100: data <= 3'b111;
            11'b01111010101: data <= 3'b111;
            11'b01111010110: data <= 3'b011;
            11'b01111010111: data <= 3'b011;
            11'b01111011000: data <= 3'b111;
            11'b01111011001: data <= 3'b111;
            11'b01111011010: data <= 3'b111;
            11'b01111011011: data <= 3'b111;
            11'b01111011100: data <= 3'b111;
            11'b01111011101: data <= 3'b110;
            11'b01111011110: data <= 3'b111;
            11'b01111011111: data <= 3'b111;
            11'b01111100000: data <= 3'b011;
            11'b01111100001: data <= 3'b011;
            11'b01111100010: data <= 3'b011;
            11'b01111100011: data <= 3'b111;
            11'b01111100100: data <= 3'b111;
            11'b01111100101: data <= 3'b111;
            11'b01111100110: data <= 3'b111;
            11'b01111100111: data <= 3'b111;
            11'b01111101000: data <= 3'b011;
            11'b01111101001: data <= 3'b111;
            11'b01111101010: data <= 3'b111;
            11'b01111101011: data <= 3'b011;
            11'b01111101100: data <= 3'b111;
            11'b01111101101: data <= 3'b111;
            11'b01111101110: data <= 3'b001;
            11'b01111101111: data <= 3'b001;
            11'b01111110000: data <= 3'b010;
            11'b01111110001: data <= 3'b010;
            11'b01111110010: data <= 3'b001;
            11'b01111110011: data <= 3'b001;
            11'b01111110100: data <= 3'b001;
            11'b01111110101: data <= 3'b001;
            11'b01111110110: data <= 3'b001;
            11'b01111110111: data <= 3'b001;
            11'b01111111000: data <= 3'b001;
            11'b01111111001: data <= 3'b001;
            11'b01111111010: data <= 3'b001;
            11'b01111111011: data <= 3'b001;
            11'b01111111100: data <= 3'b001;
            11'b01111111101: data <= 3'b001;
            11'b01111111110: data <= 3'b001;
            11'b01111111111: data <= 3'b001;
            11'b10000000000: data <= 3'b001;
            11'b10000000001: data <= 3'b001;
            11'b10000000010: data <= 3'b001;
            11'b10000000011: data <= 3'b001;
            11'b10000000100: data <= 3'b001;
            11'b10000000101: data <= 3'b001;
            11'b10000000110: data <= 3'b001;
            11'b10000000111: data <= 3'b001;
            11'b10000001000: data <= 3'b001;
            11'b10000001001: data <= 3'b001;
            11'b10000001010: data <= 3'b001;
            11'b10000001011: data <= 3'b001;
            11'b10000001100: data <= 3'b001;
            11'b10000001101: data <= 3'b000;
            11'b10000001110: data <= 3'b000;
            11'b10000001111: data <= 3'b001;
            11'b10000010000: data <= 3'b001;
            11'b10000010001: data <= 3'b001;
            11'b10000010010: data <= 3'b001;
            11'b10000010011: data <= 3'b111;
            11'b10000010100: data <= 3'b001;
            11'b10000010101: data <= 3'b011;
            11'b10000010110: data <= 3'b111;
            11'b10000010111: data <= 3'b111;
            11'b10000011000: data <= 3'b111;
            11'b10000011001: data <= 3'b001;
            11'b10000011010: data <= 3'b111;
            11'b10000011011: data <= 3'b111;
            11'b10000011100: data <= 3'b111;
            11'b10000011101: data <= 3'b111;
            11'b10000011110: data <= 3'b111;
            11'b10000011111: data <= 3'b111;
            11'b10000100000: data <= 3'b111;
            11'b10000100001: data <= 3'b111;
            11'b10000100010: data <= 3'b111;
            11'b10000100011: data <= 3'b111;
            11'b10000100100: data <= 3'b111;
            11'b10000100101: data <= 3'b111;
            11'b10000100110: data <= 3'b011;
            11'b10000100111: data <= 3'b111;
            11'b10000101000: data <= 3'b111;
            11'b10000101001: data <= 3'b011;
            11'b10000101010: data <= 3'b001;
            11'b10000101011: data <= 3'b111;
            11'b10000101100: data <= 3'b011;
            11'b10000101101: data <= 3'b001;
            11'b10000101110: data <= 3'b001;
            11'b10000101111: data <= 3'b001;
            11'b10000110000: data <= 3'b001;
            11'b10000110001: data <= 3'b000;
            11'b10000110010: data <= 3'b001;
            11'b10000110011: data <= 3'b001;
            11'b10000110100: data <= 3'b001;
            11'b10000110101: data <= 3'b001;
            11'b10000110110: data <= 3'b001;
            11'b10000110111: data <= 3'b001;
            11'b10000111000: data <= 3'b001;
            11'b10000111001: data <= 3'b001;
            11'b10000111010: data <= 3'b001;
            11'b10000111011: data <= 3'b001;
            11'b10000111100: data <= 3'b001;
            11'b10000111101: data <= 3'b001;
            11'b10000111110: data <= 3'b001;
            11'b10000111111: data <= 3'b001;
            11'b10001000000: data <= 3'b001;
            11'b10001000001: data <= 3'b001;
            11'b10001000010: data <= 3'b001;
            11'b10001000011: data <= 3'b001;
            11'b10001000100: data <= 3'b001;
            11'b10001000101: data <= 3'b001;
            11'b10001000110: data <= 3'b001;
            11'b10001000111: data <= 3'b001;
            11'b10001001000: data <= 3'b001;
            11'b10001001001: data <= 3'b001;
            11'b10001001010: data <= 3'b001;
            11'b10001001011: data <= 3'b001;
            11'b10001001100: data <= 3'b001;
            11'b10001001101: data <= 3'b001;
            11'b10001001110: data <= 3'b001;
            11'b10001001111: data <= 3'b001;
            11'b10001010000: data <= 3'b001;
            11'b10001010001: data <= 3'b001;
            11'b10001010010: data <= 3'b001;
            11'b10001010011: data <= 3'b001;
            11'b10001010100: data <= 3'b001;
            11'b10001010101: data <= 3'b001;
            11'b10001010110: data <= 3'b111;
            11'b10001010111: data <= 3'b111;
            11'b10001011000: data <= 3'b111;
            11'b10001011001: data <= 3'b001;
            11'b10001011010: data <= 3'b001;
            11'b10001011011: data <= 3'b001;
            11'b10001011100: data <= 3'b001;
            11'b10001011101: data <= 3'b001;
            11'b10001011110: data <= 3'b011;
            11'b10001011111: data <= 3'b001;
            11'b10001100000: data <= 3'b011;
            11'b10001100001: data <= 3'b001;
            11'b10001100010: data <= 3'b001;
            11'b10001100011: data <= 3'b001;
            11'b10001100100: data <= 3'b001;
            11'b10001100101: data <= 3'b001;
            11'b10001100110: data <= 3'b111;
            11'b10001100111: data <= 3'b111;
            11'b10001101000: data <= 3'b111;
            11'b10001101001: data <= 3'b001;
            11'b10001101010: data <= 3'b001;
            11'b10001101011: data <= 3'b001;
            11'b10001101100: data <= 3'b001;
            11'b10001101101: data <= 3'b001;
            11'b10001101110: data <= 3'b001;
            11'b10001101111: data <= 3'b001;
            11'b10001110000: data <= 3'b001;
            11'b10001110001: data <= 3'b001;
            11'b10001110010: data <= 3'b001;
            11'b10001110011: data <= 3'b001;
            11'b10001110100: data <= 3'b001;
            11'b10001110101: data <= 3'b001;
            11'b10001110110: data <= 3'b001;
            11'b10001110111: data <= 3'b001;
            11'b10001111000: data <= 3'b001;
            11'b10001111001: data <= 3'b001;
            11'b10001111010: data <= 3'b001;
            11'b10001111011: data <= 3'b001;
            11'b10001111100: data <= 3'b001;
            11'b10001111101: data <= 3'b001;
            11'b10001111110: data <= 3'b001;
            11'b10001111111: data <= 3'b001;
            11'b10010000000: data <= 3'b001;
            11'b10010000001: data <= 3'b001;
            11'b10010000010: data <= 3'b001;
            11'b10010000011: data <= 3'b001;
            11'b10010000100: data <= 3'b001;
            11'b10010000101: data <= 3'b001;
            11'b10010000110: data <= 3'b001;
            11'b10010000111: data <= 3'b001;
            11'b10010001000: data <= 3'b001;
            11'b10010001001: data <= 3'b001;
            11'b10010001010: data <= 3'b001;
            11'b10010001011: data <= 3'b001;
            11'b10010001100: data <= 3'b001;
            11'b10010001101: data <= 3'b001;
            11'b10010001110: data <= 3'b001;
            11'b10010001111: data <= 3'b001;
            11'b10010010000: data <= 3'b001;
            11'b10010010001: data <= 3'b001;
            11'b10010010010: data <= 3'b001;
            11'b10010010011: data <= 3'b001;
            11'b10010010100: data <= 3'b001;
            11'b10010010101: data <= 3'b001;
            11'b10010010110: data <= 3'b011;
            11'b10010010111: data <= 3'b010;
            11'b10010011000: data <= 3'b111;
            11'b10010011001: data <= 3'b111;
            11'b10010011010: data <= 3'b011;
            11'b10010011011: data <= 3'b001;
            11'b10010011100: data <= 3'b001;
            11'b10010011101: data <= 3'b001;
            11'b10010011110: data <= 3'b001;
            11'b10010011111: data <= 3'b001;
            11'b10010100000: data <= 3'b001;
            11'b10010100001: data <= 3'b001;
            11'b10010100010: data <= 3'b001;
            11'b10010100011: data <= 3'b001;
            11'b10010100100: data <= 3'b001;
            11'b10010100101: data <= 3'b111;
            11'b10010100110: data <= 3'b111;
            11'b10010100111: data <= 3'b010;
            11'b10010101000: data <= 3'b011;
            11'b10010101001: data <= 3'b001;
            11'b10010101010: data <= 3'b001;
            11'b10010101011: data <= 3'b001;
            11'b10010101100: data <= 3'b001;
            11'b10010101101: data <= 3'b001;
            11'b10010101110: data <= 3'b001;
            11'b10010101111: data <= 3'b001;
            11'b10010110000: data <= 3'b001;
            11'b10010110001: data <= 3'b001;
            11'b10010110010: data <= 3'b001;
            11'b10010110011: data <= 3'b001;
            11'b10010110100: data <= 3'b001;
            11'b10010110101: data <= 3'b001;
            11'b10010110110: data <= 3'b001;
            11'b10010110111: data <= 3'b001;
            11'b10010111000: data <= 3'b001;
            11'b10010111001: data <= 3'b001;
            11'b10010111010: data <= 3'b001;
            11'b10010111011: data <= 3'b001;
            11'b10010111100: data <= 3'b001;
            11'b10010111101: data <= 3'b001;
            11'b10010111110: data <= 3'b001;
            11'b10010111111: data <= 3'b001;
            11'b10011000000: data <= 3'b001;
            11'b10011000001: data <= 3'b001;
            11'b10011000010: data <= 3'b001;
            11'b10011000011: data <= 3'b001;
            11'b10011000100: data <= 3'b001;
            11'b10011000101: data <= 3'b001;
            11'b10011000110: data <= 3'b001;
            11'b10011000111: data <= 3'b001;
            11'b10011001000: data <= 3'b001;
            11'b10011001001: data <= 3'b001;
            11'b10011001010: data <= 3'b001;
            11'b10011001011: data <= 3'b001;
            11'b10011001100: data <= 3'b001;
            11'b10011001101: data <= 3'b001;
            11'b10011001110: data <= 3'b001;
            11'b10011001111: data <= 3'b001;
            11'b10011010000: data <= 3'b001;
            11'b10011010001: data <= 3'b001;
            11'b10011010010: data <= 3'b001;
            11'b10011010011: data <= 3'b001;
            11'b10011010100: data <= 3'b001;
            11'b10011010101: data <= 3'b001;
            11'b10011010110: data <= 3'b001;
            11'b10011010111: data <= 3'b001;
            11'b10011011000: data <= 3'b001;
            11'b10011011001: data <= 3'b111;
            11'b10011011010: data <= 3'b111;
            11'b10011011011: data <= 3'b111;
            11'b10011011100: data <= 3'b001;
            11'b10011011101: data <= 3'b111;
            11'b10011011110: data <= 3'b011;
            11'b10011011111: data <= 3'b001;
            11'b10011100000: data <= 3'b001;
            11'b10011100001: data <= 3'b111;
            11'b10011100010: data <= 3'b001;
            11'b10011100011: data <= 3'b111;
            11'b10011100100: data <= 3'b111;
            11'b10011100101: data <= 3'b111;
            11'b10011100110: data <= 3'b001;
            11'b10011100111: data <= 3'b001;
            11'b10011101000: data <= 3'b001;
            11'b10011101001: data <= 3'b001;
            11'b10011101010: data <= 3'b001;
            11'b10011101011: data <= 3'b001;
            11'b10011101100: data <= 3'b001;
            11'b10011101101: data <= 3'b001;
            11'b10011101110: data <= 3'b001;
            11'b10011101111: data <= 3'b001;
            11'b10011110000: data <= 3'b001;
            11'b10011110001: data <= 3'b001;
            11'b10011110010: data <= 3'b001;
            11'b10011110011: data <= 3'b001;
            11'b10011110100: data <= 3'b001;
            11'b10011110101: data <= 3'b001;
            11'b10011110110: data <= 3'b001;
            11'b10011110111: data <= 3'b001;
            11'b10011111000: data <= 3'b001;
            11'b10011111001: data <= 3'b001;
            11'b10011111010: data <= 3'b001;
            11'b10011111011: data <= 3'b001;
            11'b10011111100: data <= 3'b001;
            11'b10011111101: data <= 3'b001;
            11'b10011111110: data <= 3'b001;
            11'b10011111111: data <= 3'b001;
            11'b10100000000: data <= 3'b001;
            11'b10100000001: data <= 3'b001;
            11'b10100000010: data <= 3'b001;
            11'b10100000011: data <= 3'b001;
            11'b10100000100: data <= 3'b001;
            11'b10100000101: data <= 3'b001;
            11'b10100000110: data <= 3'b001;
            11'b10100000111: data <= 3'b001;
            11'b10100001000: data <= 3'b001;
            11'b10100001001: data <= 3'b001;
            11'b10100001010: data <= 3'b001;
            11'b10100001011: data <= 3'b001;
            11'b10100001100: data <= 3'b001;
            11'b10100001101: data <= 3'b001;
            11'b10100001110: data <= 3'b001;
            11'b10100001111: data <= 3'b001;
            11'b10100010000: data <= 3'b001;
            11'b10100010001: data <= 3'b001;
            11'b10100010010: data <= 3'b001;
            11'b10100010011: data <= 3'b001;
            11'b10100010100: data <= 3'b001;
            11'b10100010101: data <= 3'b001;
            11'b10100010110: data <= 3'b001;
            11'b10100010111: data <= 3'b001;
            11'b10100011000: data <= 3'b001;
            11'b10100011001: data <= 3'b001;
            11'b10100011010: data <= 3'b000;
            11'b10100011011: data <= 3'b111;
            11'b10100011100: data <= 3'b001;
            11'b10100011101: data <= 3'b001;
            11'b10100011110: data <= 3'b001;
            11'b10100011111: data <= 3'b001;
            11'b10100100000: data <= 3'b001;
            11'b10100100001: data <= 3'b001;
            11'b10100100010: data <= 3'b001;
            11'b10100100011: data <= 3'b111;
            11'b10100100100: data <= 3'b010;
            11'b10100100101: data <= 3'b001;
            11'b10100100110: data <= 3'b001;
            11'b10100100111: data <= 3'b001;
            11'b10100101000: data <= 3'b001;
            11'b10100101001: data <= 3'b001;
            11'b10100101010: data <= 3'b001;
            11'b10100101011: data <= 3'b001;
            11'b10100101100: data <= 3'b001;
            11'b10100101101: data <= 3'b001;
            11'b10100101110: data <= 3'b001;
            11'b10100101111: data <= 3'b001;
            11'b10100110000: data <= 3'b001;
            11'b10100110001: data <= 3'b001;
            11'b10100110010: data <= 3'b001;
            11'b10100110011: data <= 3'b001;
            11'b10100110100: data <= 3'b001;
            11'b10100110101: data <= 3'b001;
            11'b10100110110: data <= 3'b001;
            11'b10100110111: data <= 3'b001;
            11'b10100111000: data <= 3'b001;
            11'b10100111001: data <= 3'b001;
            11'b10100111010: data <= 3'b001;
            11'b10100111011: data <= 3'b001;
            11'b10100111100: data <= 3'b001;
            11'b10100111101: data <= 3'b001;
            11'b10100111110: data <= 3'b001;
            11'b10100111111: data <= 3'b001;
            11'b10101000000: data <= 3'b001;
            11'b10101000001: data <= 3'b001;
            11'b10101000010: data <= 3'b001;
            11'b10101000011: data <= 3'b001;
            11'b10101000100: data <= 3'b001;
            11'b10101000101: data <= 3'b001;
            11'b10101000110: data <= 3'b001;
            11'b10101000111: data <= 3'b001;
            11'b10101001000: data <= 3'b001;
            11'b10101001001: data <= 3'b001;
            11'b10101001010: data <= 3'b001;
            11'b10101001011: data <= 3'b001;
            11'b10101001100: data <= 3'b001;
            11'b10101001101: data <= 3'b001;
            11'b10101001110: data <= 3'b001;
            11'b10101001111: data <= 3'b001;
            11'b10101010000: data <= 3'b001;
            11'b10101010001: data <= 3'b001;
            11'b10101010010: data <= 3'b001;
            11'b10101010011: data <= 3'b001;
            11'b10101010100: data <= 3'b001;
            11'b10101010101: data <= 3'b001;
            11'b10101010110: data <= 3'b001;
            11'b10101010111: data <= 3'b001;
            11'b10101011000: data <= 3'b001;
            11'b10101011001: data <= 3'b001;
            11'b10101011010: data <= 3'b001;
            11'b10101011011: data <= 3'b001;
            11'b10101011100: data <= 3'b001;
            11'b10101011101: data <= 3'b001;
            11'b10101011110: data <= 3'b001;
            11'b10101011111: data <= 3'b001;
            11'b10101100000: data <= 3'b001;
            11'b10101100001: data <= 3'b001;
            11'b10101100010: data <= 3'b001;
            11'b10101100011: data <= 3'b001;
            11'b10101100100: data <= 3'b001;
            11'b10101100101: data <= 3'b001;
            11'b10101100110: data <= 3'b001;
            11'b10101100111: data <= 3'b001;
            11'b10101101000: data <= 3'b001;
            11'b10101101001: data <= 3'b001;
            11'b10101101010: data <= 3'b001;
            11'b10101101011: data <= 3'b001;
            11'b10101101100: data <= 3'b001;
            11'b10101101101: data <= 3'b001;
            11'b10101101110: data <= 3'b001;
            11'b10101101111: data <= 3'b001;
            11'b10101110000: data <= 3'b001;
            11'b10101110001: data <= 3'b001;
            11'b10101110010: data <= 3'b001;
            11'b10101110011: data <= 3'b001;
            11'b10101110100: data <= 3'b001;
            11'b10101110101: data <= 3'b001;
            11'b10101110110: data <= 3'b001;
            11'b10101110111: data <= 3'b001;
            11'b10101111000: data <= 3'b001;
            11'b10101111001: data <= 3'b001;
            11'b10101111010: data <= 3'b001;
            11'b10101111011: data <= 3'b001;
            11'b10101111100: data <= 3'b001;
            11'b10101111101: data <= 3'b001;
            11'b10101111110: data <= 3'b001;
            11'b10101111111: data <= 3'b001;
            11'b10110000000: data <= 3'b001;
            11'b10110000001: data <= 3'b001;
            11'b10110000010: data <= 3'b001;
            11'b10110000011: data <= 3'b001;
            11'b10110000100: data <= 3'b001;
            11'b10110000101: data <= 3'b001;
            11'b10110000110: data <= 3'b001;
            11'b10110000111: data <= 3'b001;
            11'b10110001000: data <= 3'b001;
            11'b10110001001: data <= 3'b001;
            11'b10110001010: data <= 3'b001;
            11'b10110001011: data <= 3'b001;
            11'b10110001100: data <= 3'b001;
            11'b10110001101: data <= 3'b001;
            11'b10110001110: data <= 3'b001;
            11'b10110001111: data <= 3'b001;
            11'b10110010000: data <= 3'b001;
            11'b10110010001: data <= 3'b001;
            11'b10110010010: data <= 3'b001;
            11'b10110010011: data <= 3'b001;
            11'b10110010100: data <= 3'b001;
            11'b10110010101: data <= 3'b001;
            11'b10110010110: data <= 3'b001;
            11'b10110010111: data <= 3'b001;
            11'b10110011000: data <= 3'b001;
            11'b10110011001: data <= 3'b001;
            11'b10110011010: data <= 3'b001;
            11'b10110011011: data <= 3'b001;
            11'b10110011100: data <= 3'b001;
            11'b10110011101: data <= 3'b001;
            11'b10110011110: data <= 3'b001;
            11'b10110011111: data <= 3'b001;
            11'b10110100000: data <= 3'b001;
            11'b10110100001: data <= 3'b001;
            11'b10110100010: data <= 3'b001;
            11'b10110100011: data <= 3'b001;
            11'b10110100100: data <= 3'b001;
            11'b10110100101: data <= 3'b001;
            11'b10110100110: data <= 3'b001;
            11'b10110100111: data <= 3'b001;
            11'b10110101000: data <= 3'b001;
            11'b10110101001: data <= 3'b001;
            11'b10110101010: data <= 3'b001;
            11'b10110101011: data <= 3'b001;
            11'b10110101100: data <= 3'b001;
            11'b10110101101: data <= 3'b001;
            11'b10110101110: data <= 3'b001;
            11'b10110101111: data <= 3'b001;
            11'b10110110000: data <= 3'b001;
            11'b10110110001: data <= 3'b001;
            11'b10110110010: data <= 3'b001;
            11'b10110110011: data <= 3'b001;
            11'b10110110100: data <= 3'b001;
            11'b10110110101: data <= 3'b001;
            11'b10110110110: data <= 3'b001;
            11'b10110110111: data <= 3'b001;
            11'b10110111000: data <= 3'b001;
            11'b10110111001: data <= 3'b001;
            11'b10110111010: data <= 3'b001;
            11'b10110111011: data <= 3'b001;
            11'b10110111100: data <= 3'b001;
            11'b10110111101: data <= 3'b001;
            11'b10110111110: data <= 3'b001;
            11'b10110111111: data <= 3'b001;
            11'b10111000000: data <= 3'b001;
            11'b10111000001: data <= 3'b001;
            11'b10111000010: data <= 3'b001;
            11'b10111000011: data <= 3'b001;
            11'b10111000100: data <= 3'b001;
            11'b10111000101: data <= 3'b001;
            11'b10111000110: data <= 3'b001;
            11'b10111000111: data <= 3'b001;
            11'b10111001000: data <= 3'b001;
            11'b10111001001: data <= 3'b001;
            11'b10111001010: data <= 3'b001;
            11'b10111001011: data <= 3'b001;
            11'b10111001100: data <= 3'b001;
            11'b10111001101: data <= 3'b001;
            11'b10111001110: data <= 3'b001;
            11'b10111001111: data <= 3'b001;
            11'b10111010000: data <= 3'b001;
            11'b10111010001: data <= 3'b001;
            11'b10111010010: data <= 3'b001;
            11'b10111010011: data <= 3'b001;
            11'b10111010100: data <= 3'b001;
            11'b10111010101: data <= 3'b001;
            11'b10111010110: data <= 3'b001;
            11'b10111010111: data <= 3'b001;
            11'b10111011000: data <= 3'b001;
            11'b10111011001: data <= 3'b001;
            11'b10111011010: data <= 3'b001;
            11'b10111011011: data <= 3'b001;
            11'b10111011100: data <= 3'b001;
            11'b10111011101: data <= 3'b001;
            11'b10111011110: data <= 3'b001;
            11'b10111011111: data <= 3'b001;
            11'b10111100000: data <= 3'b001;
            11'b10111100001: data <= 3'b001;
            11'b10111100010: data <= 3'b001;
            11'b10111100011: data <= 3'b001;
            11'b10111100100: data <= 3'b001;
            11'b10111100101: data <= 3'b001;
            11'b10111100110: data <= 3'b001;
            11'b10111100111: data <= 3'b001;
            11'b10111101000: data <= 3'b001;
            11'b10111101001: data <= 3'b001;
            11'b10111101010: data <= 3'b001;
            11'b10111101011: data <= 3'b001;
            11'b10111101100: data <= 3'b001;
            11'b10111101101: data <= 3'b001;
            11'b10111101110: data <= 3'b001;
            11'b10111101111: data <= 3'b001;
            11'b10111110000: data <= 3'b001;
            11'b10111110001: data <= 3'b001;
            11'b10111110010: data <= 3'b001;
            11'b10111110011: data <= 3'b001;
            11'b10111110100: data <= 3'b001;
            11'b10111110101: data <= 3'b001;
            11'b10111110110: data <= 3'b001;
            11'b10111110111: data <= 3'b001;
            11'b10111111000: data <= 3'b001;
            11'b10111111001: data <= 3'b001;
            11'b10111111010: data <= 3'b001;
            11'b10111111011: data <= 3'b001;
            11'b10111111100: data <= 3'b001;
            11'b10111111101: data <= 3'b001;
            11'b10111111110: data <= 3'b001;
            11'b10111111111: data <= 3'b001;
            11'b11000000000: data <= 3'b001;
            11'b11000000001: data <= 3'b001;
            11'b11000000010: data <= 3'b001;
            11'b11000000011: data <= 3'b001;
            11'b11000000100: data <= 3'b001;
            11'b11000000101: data <= 3'b001;
            11'b11000000110: data <= 3'b001;
            11'b11000000111: data <= 3'b001;
            11'b11000001000: data <= 3'b001;
            11'b11000001001: data <= 3'b001;
            11'b11000001010: data <= 3'b001;
            11'b11000001011: data <= 3'b001;
            11'b11000001100: data <= 3'b001;
            11'b11000001101: data <= 3'b001;
            11'b11000001110: data <= 3'b001;
            11'b11000001111: data <= 3'b001;
            11'b11000010000: data <= 3'b001;
            11'b11000010001: data <= 3'b001;
            11'b11000010010: data <= 3'b001;
            11'b11000010011: data <= 3'b001;
            11'b11000010100: data <= 3'b001;
            11'b11000010101: data <= 3'b001;
            11'b11000010110: data <= 3'b001;
            11'b11000010111: data <= 3'b001;
            11'b11000011000: data <= 3'b001;
            11'b11000011001: data <= 3'b001;
            11'b11000011010: data <= 3'b001;
            11'b11000011011: data <= 3'b001;
            11'b11000011100: data <= 3'b001;
            11'b11000011101: data <= 3'b001;
            11'b11000011110: data <= 3'b001;
            11'b11000011111: data <= 3'b001;
            11'b11000100000: data <= 3'b001;
            11'b11000100001: data <= 3'b001;
            11'b11000100010: data <= 3'b001;
            11'b11000100011: data <= 3'b001;
            11'b11000100100: data <= 3'b001;
            11'b11000100101: data <= 3'b001;
            11'b11000100110: data <= 3'b001;
            11'b11000100111: data <= 3'b001;
            11'b11000101000: data <= 3'b001;
            11'b11000101001: data <= 3'b001;
            11'b11000101010: data <= 3'b001;
            11'b11000101011: data <= 3'b001;
            11'b11000101100: data <= 3'b001;
            11'b11000101101: data <= 3'b001;
            11'b11000101110: data <= 3'b001;
            11'b11000101111: data <= 3'b001;
            11'b11000110000: data <= 3'b001;
            11'b11000110001: data <= 3'b001;
            11'b11000110010: data <= 3'b001;
            11'b11000110011: data <= 3'b001;
            11'b11000110100: data <= 3'b001;
            11'b11000110101: data <= 3'b001;
            11'b11000110110: data <= 3'b001;
            11'b11000110111: data <= 3'b001;
            11'b11000111000: data <= 3'b001;
            11'b11000111001: data <= 3'b001;
            11'b11000111010: data <= 3'b001;
            11'b11000111011: data <= 3'b001;
            11'b11000111100: data <= 3'b001;
            11'b11000111101: data <= 3'b001;
            11'b11000111110: data <= 3'b001;
            11'b11000111111: data <= 3'b001;
            11'b11001000000: data <= 3'b001;
            11'b11001000001: data <= 3'b001;
            11'b11001000010: data <= 3'b001;
            11'b11001000011: data <= 3'b001;
            11'b11001000100: data <= 3'b001;
            11'b11001000101: data <= 3'b001;
            11'b11001000110: data <= 3'b001;
            11'b11001000111: data <= 3'b001;
            11'b11001001000: data <= 3'b001;
            11'b11001001001: data <= 3'b001;
            11'b11001001010: data <= 3'b001;
            11'b11001001011: data <= 3'b001;
            11'b11001001100: data <= 3'b001;
            11'b11001001101: data <= 3'b001;
            11'b11001001110: data <= 3'b001;
            11'b11001001111: data <= 3'b001;
            11'b11001010000: data <= 3'b001;
            11'b11001010001: data <= 3'b001;
            11'b11001010010: data <= 3'b001;
            11'b11001010011: data <= 3'b001;
            11'b11001010100: data <= 3'b001;
            11'b11001010101: data <= 3'b001;
            11'b11001010110: data <= 3'b001;
            11'b11001010111: data <= 3'b001;
            11'b11001011000: data <= 3'b001;
            11'b11001011001: data <= 3'b001;
            11'b11001011010: data <= 3'b001;
            11'b11001011011: data <= 3'b001;
            11'b11001011100: data <= 3'b001;
            11'b11001011101: data <= 3'b001;
            11'b11001011110: data <= 3'b001;
            11'b11001011111: data <= 3'b001;
            11'b11001100000: data <= 3'b001;
            11'b11001100001: data <= 3'b001;
            11'b11001100010: data <= 3'b001;
            11'b11001100011: data <= 3'b001;
            11'b11001100100: data <= 3'b001;
            11'b11001100101: data <= 3'b001;
            11'b11001100110: data <= 3'b001;
            11'b11001100111: data <= 3'b001;
            11'b11001101000: data <= 3'b001;
            11'b11001101001: data <= 3'b001;
            11'b11001101010: data <= 3'b001;
            11'b11001101011: data <= 3'b001;
            11'b11001101100: data <= 3'b001;
            11'b11001101101: data <= 3'b001;
            11'b11001101110: data <= 3'b001;
            11'b11001101111: data <= 3'b001;
            11'b11001110000: data <= 3'b001;
            11'b11001110001: data <= 3'b001;
            11'b11001110010: data <= 3'b001;
            11'b11001110011: data <= 3'b001;
            11'b11001110100: data <= 3'b001;
            11'b11001110101: data <= 3'b001;
            11'b11001110110: data <= 3'b001;
            11'b11001110111: data <= 3'b001;
            11'b11001111000: data <= 3'b001;
            11'b11001111001: data <= 3'b001;
            11'b11001111010: data <= 3'b001;
            11'b11001111011: data <= 3'b001;
            11'b11001111100: data <= 3'b001;
            11'b11001111101: data <= 3'b001;
            11'b11001111110: data <= 3'b001;
            11'b11001111111: data <= 3'b001;
            11'b11010000000: data <= 3'b001;
            11'b11010000001: data <= 3'b001;
            11'b11010000010: data <= 3'b001;
            11'b11010000011: data <= 3'b001;
            11'b11010000100: data <= 3'b001;
            11'b11010000101: data <= 3'b001;
            11'b11010000110: data <= 3'b001;
            11'b11010000111: data <= 3'b001;
            11'b11010001000: data <= 3'b001;
            11'b11010001001: data <= 3'b001;
            11'b11010001010: data <= 3'b001;
            11'b11010001011: data <= 3'b001;
            11'b11010001100: data <= 3'b001;
            11'b11010001101: data <= 3'b001;
            11'b11010001110: data <= 3'b001;
            11'b11010001111: data <= 3'b001;
            11'b11010010000: data <= 3'b001;
            11'b11010010001: data <= 3'b001;
            11'b11010010010: data <= 3'b001;
            11'b11010010011: data <= 3'b001;
            11'b11010010100: data <= 3'b001;
            11'b11010010101: data <= 3'b001;
            11'b11010010110: data <= 3'b001;
            11'b11010010111: data <= 3'b001;
            11'b11010011000: data <= 3'b001;
            11'b11010011001: data <= 3'b001;
            11'b11010011010: data <= 3'b001;
            11'b11010011011: data <= 3'b001;
            11'b11010011100: data <= 3'b001;
            11'b11010011101: data <= 3'b001;
            11'b11010011110: data <= 3'b001;
            11'b11010011111: data <= 3'b001;
            11'b11010100000: data <= 3'b001;
            11'b11010100001: data <= 3'b001;
            11'b11010100010: data <= 3'b001;
            11'b11010100011: data <= 3'b001;
            11'b11010100100: data <= 3'b001;
            11'b11010100101: data <= 3'b001;
            11'b11010100110: data <= 3'b001;
            11'b11010100111: data <= 3'b001;
            11'b11010101000: data <= 3'b001;
            11'b11010101001: data <= 3'b001;
            11'b11010101010: data <= 3'b001;
            11'b11010101011: data <= 3'b001;
            11'b11010101100: data <= 3'b001;
            11'b11010101101: data <= 3'b001;
            11'b11010101110: data <= 3'b001;
            11'b11010101111: data <= 3'b001;
            11'b11010110000: data <= 3'b001;
            11'b11010110001: data <= 3'b001;
            11'b11010110010: data <= 3'b001;
            11'b11010110011: data <= 3'b001;
            11'b11010110100: data <= 3'b001;
            11'b11010110101: data <= 3'b001;
            11'b11010110110: data <= 3'b001;
            11'b11010110111: data <= 3'b001;
            11'b11010111000: data <= 3'b001;
            11'b11010111001: data <= 3'b001;
            11'b11010111010: data <= 3'b001;
            11'b11010111011: data <= 3'b001;
            11'b11010111100: data <= 3'b001;
            11'b11010111101: data <= 3'b001;
            11'b11010111110: data <= 3'b001;
            11'b11010111111: data <= 3'b001;
            11'b11011000000: data <= 3'b001;
            11'b11011000001: data <= 3'b001;
            11'b11011000010: data <= 3'b001;
            11'b11011000011: data <= 3'b001;
            11'b11011000100: data <= 3'b001;
            11'b11011000101: data <= 3'b001;
            11'b11011000110: data <= 3'b001;
            11'b11011000111: data <= 3'b001;
            11'b11011001000: data <= 3'b001;
            11'b11011001001: data <= 3'b001;
            11'b11011001010: data <= 3'b001;
            11'b11011001011: data <= 3'b001;
            11'b11011001100: data <= 3'b001;
            11'b11011001101: data <= 3'b001;
            11'b11011001110: data <= 3'b001;
            11'b11011001111: data <= 3'b001;
            11'b11011010000: data <= 3'b001;
            11'b11011010001: data <= 3'b001;
            11'b11011010010: data <= 3'b001;
            11'b11011010011: data <= 3'b001;
            11'b11011010100: data <= 3'b001;
            11'b11011010101: data <= 3'b001;
            11'b11011010110: data <= 3'b001;
            11'b11011010111: data <= 3'b001;
            11'b11011011000: data <= 3'b001;
            11'b11011011001: data <= 3'b001;
            11'b11011011010: data <= 3'b001;
            11'b11011011011: data <= 3'b001;
            11'b11011011100: data <= 3'b001;
            11'b11011011101: data <= 3'b001;
            11'b11011011110: data <= 3'b001;
            11'b11011011111: data <= 3'b001;
            11'b11011100000: data <= 3'b001;
            11'b11011100001: data <= 3'b001;
            11'b11011100010: data <= 3'b001;
            11'b11011100011: data <= 3'b001;
            11'b11011100100: data <= 3'b001;
            11'b11011100101: data <= 3'b001;
            11'b11011100110: data <= 3'b001;
            11'b11011100111: data <= 3'b001;
            11'b11011101000: data <= 3'b001;
            11'b11011101001: data <= 3'b001;
            11'b11011101010: data <= 3'b001;
            11'b11011101011: data <= 3'b001;
            11'b11011101100: data <= 3'b001;
            11'b11011101101: data <= 3'b001;
            11'b11011101110: data <= 3'b001;
            11'b11011101111: data <= 3'b001;
            11'b11011110000: data <= 3'b001;
            11'b11011110001: data <= 3'b001;
            11'b11011110010: data <= 3'b001;
            11'b11011110011: data <= 3'b001;
            11'b11011110100: data <= 3'b001;
            11'b11011110101: data <= 3'b001;
            11'b11011110110: data <= 3'b001;
            11'b11011110111: data <= 3'b001;
            11'b11011111000: data <= 3'b001;
            11'b11011111001: data <= 3'b001;
            11'b11011111010: data <= 3'b001;
            11'b11011111011: data <= 3'b001;
            11'b11011111100: data <= 3'b001;
            11'b11011111101: data <= 3'b001;
            11'b11011111110: data <= 3'b001;
            11'b11011111111: data <= 3'b001;
            11'b11100000000: data <= 3'b001;
            11'b11100000001: data <= 3'b001;
            11'b11100000010: data <= 3'b001;
            11'b11100000011: data <= 3'b001;
            11'b11100000100: data <= 3'b001;
            11'b11100000101: data <= 3'b001;
            11'b11100000110: data <= 3'b001;
            11'b11100000111: data <= 3'b001;
            11'b11100001000: data <= 3'b001;
            11'b11100001001: data <= 3'b001;
            11'b11100001010: data <= 3'b001;
            11'b11100001011: data <= 3'b001;
            11'b11100001100: data <= 3'b001;
            11'b11100001101: data <= 3'b001;
            11'b11100001110: data <= 3'b001;
            11'b11100001111: data <= 3'b001;
            11'b11100010000: data <= 3'b001;
            11'b11100010001: data <= 3'b001;
            11'b11100010010: data <= 3'b001;
            11'b11100010011: data <= 3'b001;
            11'b11100010100: data <= 3'b001;
            11'b11100010101: data <= 3'b001;
            11'b11100010110: data <= 3'b001;
            11'b11100010111: data <= 3'b001;
            11'b11100011000: data <= 3'b001;
            11'b11100011001: data <= 3'b001;
            11'b11100011010: data <= 3'b001;
            11'b11100011011: data <= 3'b001;
            11'b11100011100: data <= 3'b001;
            11'b11100011101: data <= 3'b001;
            11'b11100011110: data <= 3'b001;
            11'b11100011111: data <= 3'b001;
            11'b11100100000: data <= 3'b001;
            11'b11100100001: data <= 3'b001;
            11'b11100100010: data <= 3'b001;
            11'b11100100011: data <= 3'b001;
            11'b11100100100: data <= 3'b001;
            11'b11100100101: data <= 3'b001;
            11'b11100100110: data <= 3'b001;
            11'b11100100111: data <= 3'b001;
            11'b11100101000: data <= 3'b001;
            11'b11100101001: data <= 3'b001;
            11'b11100101010: data <= 3'b001;
            11'b11100101011: data <= 3'b001;
            11'b11100101100: data <= 3'b001;
            11'b11100101101: data <= 3'b001;
            11'b11100101110: data <= 3'b001;
            11'b11100101111: data <= 3'b001;
            11'b11100110000: data <= 3'b001;
            11'b11100110001: data <= 3'b001;
            11'b11100110010: data <= 3'b001;
            11'b11100110011: data <= 3'b001;
            11'b11100110100: data <= 3'b001;
            11'b11100110101: data <= 3'b001;
            11'b11100110110: data <= 3'b001;
            11'b11100110111: data <= 3'b001;
            11'b11100111000: data <= 3'b001;
            11'b11100111001: data <= 3'b001;
            11'b11100111010: data <= 3'b001;
            11'b11100111011: data <= 3'b001;
            11'b11100111100: data <= 3'b001;
            11'b11100111101: data <= 3'b001;
            11'b11100111110: data <= 3'b001;
            11'b11100111111: data <= 3'b001;
            11'b11101000000: data <= 3'b001;
            11'b11101000001: data <= 3'b001;
            11'b11101000010: data <= 3'b001;
            11'b11101000011: data <= 3'b001;
            11'b11101000100: data <= 3'b001;
            11'b11101000101: data <= 3'b001;
            11'b11101000110: data <= 3'b001;
            11'b11101000111: data <= 3'b001;
            11'b11101001000: data <= 3'b001;
            11'b11101001001: data <= 3'b001;
            11'b11101001010: data <= 3'b001;
            11'b11101001011: data <= 3'b001;
            11'b11101001100: data <= 3'b001;
            11'b11101001101: data <= 3'b001;
            11'b11101001110: data <= 3'b001;
            11'b11101001111: data <= 3'b001;
            11'b11101010000: data <= 3'b001;
            11'b11101010001: data <= 3'b001;
            11'b11101010010: data <= 3'b001;
            11'b11101010011: data <= 3'b001;
            11'b11101010100: data <= 3'b001;
            11'b11101010101: data <= 3'b001;
            11'b11101010110: data <= 3'b001;
            11'b11101010111: data <= 3'b001;
            11'b11101011000: data <= 3'b001;
            11'b11101011001: data <= 3'b001;
            11'b11101011010: data <= 3'b001;
            11'b11101011011: data <= 3'b001;
            11'b11101011100: data <= 3'b001;
            11'b11101011101: data <= 3'b001;
            11'b11101011110: data <= 3'b001;
            11'b11101011111: data <= 3'b001;
            11'b11101100000: data <= 3'b001;
            11'b11101100001: data <= 3'b001;
            11'b11101100010: data <= 3'b001;
            11'b11101100011: data <= 3'b001;
            11'b11101100100: data <= 3'b001;
            11'b11101100101: data <= 3'b001;
            11'b11101100110: data <= 3'b001;
            11'b11101100111: data <= 3'b001;
            11'b11101101000: data <= 3'b001;
            11'b11101101001: data <= 3'b001;
            11'b11101101010: data <= 3'b001;
            11'b11101101011: data <= 3'b001;
            11'b11101101100: data <= 3'b001;
            11'b11101101101: data <= 3'b001;
            11'b11101101110: data <= 3'b001;
            11'b11101101111: data <= 3'b001;
            11'b11101110000: data <= 3'b001;
            11'b11101110001: data <= 3'b001;
            11'b11101110010: data <= 3'b001;
            11'b11101110011: data <= 3'b001;
            11'b11101110100: data <= 3'b001;
            11'b11101110101: data <= 3'b001;
            11'b11101110110: data <= 3'b001;
            11'b11101110111: data <= 3'b001;
            11'b11101111000: data <= 3'b001;
            11'b11101111001: data <= 3'b001;
            11'b11101111010: data <= 3'b001;
            11'b11101111011: data <= 3'b001;
            11'b11101111100: data <= 3'b001;
            11'b11101111101: data <= 3'b001;
            11'b11101111110: data <= 3'b001;
            11'b11101111111: data <= 3'b001;
            11'b11110000000: data <= 3'b001;
            11'b11110000001: data <= 3'b001;
            11'b11110000010: data <= 3'b001;
            11'b11110000011: data <= 3'b001;
            11'b11110000100: data <= 3'b001;
            11'b11110000101: data <= 3'b001;
            11'b11110000110: data <= 3'b001;
            11'b11110000111: data <= 3'b001;
            11'b11110001000: data <= 3'b001;
            11'b11110001001: data <= 3'b001;
            11'b11110001010: data <= 3'b001;
            11'b11110001011: data <= 3'b001;
            11'b11110001100: data <= 3'b001;
            11'b11110001101: data <= 3'b001;
            11'b11110001110: data <= 3'b001;
            11'b11110001111: data <= 3'b001;
            11'b11110010000: data <= 3'b001;
            11'b11110010001: data <= 3'b001;
            11'b11110010010: data <= 3'b001;
            11'b11110010011: data <= 3'b001;
            11'b11110010100: data <= 3'b001;
            11'b11110010101: data <= 3'b001;
            11'b11110010110: data <= 3'b001;
            11'b11110010111: data <= 3'b001;
            11'b11110011000: data <= 3'b001;
            11'b11110011001: data <= 3'b001;
            11'b11110011010: data <= 3'b001;
            11'b11110011011: data <= 3'b001;
            11'b11110011100: data <= 3'b001;
            11'b11110011101: data <= 3'b001;
            11'b11110011110: data <= 3'b001;
            11'b11110011111: data <= 3'b001;
            11'b11110100000: data <= 3'b001;
            11'b11110100001: data <= 3'b001;
            11'b11110100010: data <= 3'b001;
            11'b11110100011: data <= 3'b001;
            11'b11110100100: data <= 3'b001;
            11'b11110100101: data <= 3'b001;
            11'b11110100110: data <= 3'b001;
            11'b11110100111: data <= 3'b001;
            11'b11110101000: data <= 3'b001;
            11'b11110101001: data <= 3'b001;
            11'b11110101010: data <= 3'b001;
            11'b11110101011: data <= 3'b001;
            11'b11110101100: data <= 3'b001;
            11'b11110101101: data <= 3'b001;
            11'b11110101110: data <= 3'b001;
            11'b11110101111: data <= 3'b001;
            11'b11110110000: data <= 3'b001;
            11'b11110110001: data <= 3'b001;
            11'b11110110010: data <= 3'b001;
            11'b11110110011: data <= 3'b001;
            11'b11110110100: data <= 3'b001;
            11'b11110110101: data <= 3'b001;
            11'b11110110110: data <= 3'b001;
            11'b11110110111: data <= 3'b001;
            11'b11110111000: data <= 3'b001;
            11'b11110111001: data <= 3'b001;
            11'b11110111010: data <= 3'b001;
            11'b11110111011: data <= 3'b001;
            11'b11110111100: data <= 3'b001;
            11'b11110111101: data <= 3'b001;
            11'b11110111110: data <= 3'b001;
            11'b11110111111: data <= 3'b001;
            11'b11111000000: data <= 3'b001;
            11'b11111000001: data <= 3'b001;
            11'b11111000010: data <= 3'b001;
            11'b11111000011: data <= 3'b001;
            11'b11111000100: data <= 3'b001;
            11'b11111000101: data <= 3'b001;
            11'b11111000110: data <= 3'b001;
            11'b11111000111: data <= 3'b001;
            11'b11111001000: data <= 3'b001;
            11'b11111001001: data <= 3'b001;
            11'b11111001010: data <= 3'b001;
            11'b11111001011: data <= 3'b001;
            11'b11111001100: data <= 3'b001;
            11'b11111001101: data <= 3'b001;
            11'b11111001110: data <= 3'b001;
            11'b11111001111: data <= 3'b001;
            11'b11111010000: data <= 3'b001;
            11'b11111010001: data <= 3'b001;
            11'b11111010010: data <= 3'b001;
            11'b11111010011: data <= 3'b001;
            11'b11111010100: data <= 3'b001;
            11'b11111010101: data <= 3'b001;
            11'b11111010110: data <= 3'b001;
            11'b11111010111: data <= 3'b001;
            11'b11111011000: data <= 3'b001;
            11'b11111011001: data <= 3'b001;
            11'b11111011010: data <= 3'b001;
            11'b11111011011: data <= 3'b001;
            11'b11111011100: data <= 3'b001;
            11'b11111011101: data <= 3'b001;
            11'b11111011110: data <= 3'b001;
            11'b11111011111: data <= 3'b001;
            11'b11111100000: data <= 3'b001;
            11'b11111100001: data <= 3'b001;
            11'b11111100010: data <= 3'b001;
            11'b11111100011: data <= 3'b001;
            11'b11111100100: data <= 3'b001;
            11'b11111100101: data <= 3'b001;
            11'b11111100110: data <= 3'b001;
            11'b11111100111: data <= 3'b001;
            11'b11111101000: data <= 3'b001;
            11'b11111101001: data <= 3'b001;
            11'b11111101010: data <= 3'b001;
            11'b11111101011: data <= 3'b001;
            11'b11111101100: data <= 3'b001;
            11'b11111101101: data <= 3'b001;
            11'b11111101110: data <= 3'b001;
            11'b11111101111: data <= 3'b001;
            11'b11111110000: data <= 3'b001;
            11'b11111110001: data <= 3'b001;
            11'b11111110010: data <= 3'b001;
            11'b11111110011: data <= 3'b001;
            11'b11111110100: data <= 3'b001;
            11'b11111110101: data <= 3'b001;
            11'b11111110110: data <= 3'b001;
            11'b11111110111: data <= 3'b001;
            11'b11111111000: data <= 3'b001;
            11'b11111111001: data <= 3'b001;
            11'b11111111010: data <= 3'b001;
            11'b11111111011: data <= 3'b001;
            11'b11111111100: data <= 3'b001;
            11'b11111111101: data <= 3'b001;
            11'b11111111110: data <= 3'b001;
            11'b11111111111: data <= 3'b001;
            default: data = 3'b000;
        endcase
    end
endmodule
